magic
tech scmos
timestamp 1678804997
<< nwell >>
rect 58 42 127 73
rect 58 35 85 42
<< polysilicon >>
rect 95 59 97 61
rect 103 59 105 61
rect 111 59 113 61
rect 70 51 72 53
rect 70 41 72 43
rect 95 41 97 43
rect 70 39 97 41
rect 70 33 72 39
rect 62 29 72 33
rect 70 27 72 29
rect 98 28 100 33
rect 103 32 105 43
rect 103 30 107 32
rect 98 26 103 28
rect 101 24 103 26
rect 105 24 107 30
rect 111 27 113 43
rect 109 25 113 27
rect 109 24 111 25
rect 70 21 72 23
rect 101 10 103 12
rect 105 -6 107 12
rect 109 -6 111 12
<< ndiffusion >>
rect 64 23 65 27
rect 69 23 70 27
rect 72 23 73 27
rect 77 23 78 27
rect 95 18 101 24
rect 95 14 96 18
rect 100 14 101 18
rect 95 12 101 14
rect 103 12 105 24
rect 107 12 109 24
rect 111 18 118 24
rect 111 14 112 18
rect 116 14 118 18
rect 111 12 118 14
<< pdiffusion >>
rect 90 58 95 59
rect 94 54 95 58
rect 64 47 65 51
rect 69 47 70 51
rect 64 43 70 47
rect 72 47 73 51
rect 77 47 78 51
rect 72 43 78 47
rect 90 43 95 54
rect 97 58 103 59
rect 97 54 98 58
rect 102 54 103 58
rect 97 43 103 54
rect 105 49 111 59
rect 105 45 106 49
rect 110 45 111 49
rect 105 43 111 45
rect 113 58 118 59
rect 113 54 114 58
rect 113 43 118 54
<< metal1 >>
rect 61 71 127 73
rect 61 67 65 71
rect 69 67 90 71
rect 94 67 114 71
rect 118 67 127 71
rect 61 65 127 67
rect 65 51 69 65
rect 90 58 94 65
rect 102 54 114 58
rect 73 33 77 47
rect 106 40 110 45
rect 106 36 124 40
rect 120 33 124 36
rect 73 29 94 33
rect 73 27 77 29
rect 120 28 127 33
rect 65 9 69 23
rect 120 18 124 28
rect 116 14 124 18
rect 96 9 100 14
rect 61 8 127 9
rect 61 4 65 8
rect 69 7 127 8
rect 69 4 96 7
rect 61 3 96 4
rect 100 3 127 7
rect 61 1 127 3
<< ntransistor >>
rect 70 23 72 27
rect 101 12 103 24
rect 105 12 107 24
rect 109 12 111 24
<< ptransistor >>
rect 70 43 72 51
rect 95 43 97 59
rect 103 43 105 59
rect 111 43 113 59
<< polycontact >>
rect 58 29 62 33
rect 94 29 98 33
rect 101 -6 105 -2
rect 111 -6 115 -2
<< ndcontact >>
rect 65 23 69 27
rect 73 23 77 27
rect 96 14 100 18
rect 112 14 116 18
<< pdcontact >>
rect 90 54 94 58
rect 65 47 69 51
rect 73 47 77 51
rect 98 54 102 58
rect 106 45 110 49
rect 114 54 118 58
<< psubstratepcontact >>
rect 65 4 69 8
rect 96 3 100 7
<< nsubstratencontact >>
rect 65 67 69 71
rect 90 67 94 71
rect 114 67 118 71
<< labels >>
rlabel polycontact 58 29 62 33 7 sleep
rlabel metal1 124 28 127 33 3 out
rlabel polycontact 101 -6 105 -2 7 a
rlabel polycontact 111 -6 115 -2 3 b
rlabel metal1 61 1 127 9 5 vss
rlabel nwell 61 65 127 73 1 vdd
<< end >>
