* SPICE3 file created from nand_stt.ext - technology: scmos

.option scale=1u

M1000 a_107_12# a a_103_12# Gnd nfet w=12 l=2
+  ad=24 pd=28 as=24 ps=28
M1001 out a a_97_43# vdd pfet w=16 l=2
+  ad=96 pd=44 as=176 ps=86
M1002 a_103_12# a_72_23# vss Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=56
M1003 a_72_23# sleep vss Gnd nfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1004 a_72_23# sleep vdd vdd pfet w=8 l=2
+  ad=48 pd=28 as=128 ps=70
M1005 a_97_43# b out vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out b a_107_12# Gnd nfet w=12 l=2
+  ad=84 pd=38 as=0 ps=0
M1007 a_97_43# sleep vdd vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
C0 sleep vdd 6.99fF
C1 vss Gnd 25.00fF
C2 out Gnd 8.60fF
C3 a_72_23# Gnd 9.94fF
C4 b Gnd 10.79fF
C5 a Gnd 10.79fF
C6 sleep Gnd 9.75fF
