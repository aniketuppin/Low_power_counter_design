magic
tech scmos
timestamp 1679322495
<< nwell >>
rect -146 203 -119 241
rect -101 162 -45 199
rect -36 164 -10 205
rect -141 120 -114 161
rect 43 140 112 171
rect 144 140 213 171
rect 43 133 70 140
rect 144 133 171 140
rect 0 86 27 127
rect -103 58 -76 61
rect -30 58 -3 61
rect -103 27 -3 58
rect 46 48 115 79
rect 144 48 213 79
rect 46 41 73 48
rect 144 41 171 48
rect -103 20 -76 27
rect -30 20 -3 27
<< polysilicon >>
rect -134 221 57 223
rect -134 219 -132 221
rect -47 211 -41 212
rect -134 201 -132 211
rect -142 197 -132 201
rect -47 207 -45 211
rect -47 206 -41 207
rect -134 195 -132 197
rect -47 193 -45 206
rect -66 191 -45 193
rect -134 189 -132 191
rect -112 189 -88 191
rect -134 187 -110 189
rect -90 187 -88 189
rect -82 187 -80 189
rect -74 187 -72 189
rect -66 187 -64 191
rect -58 187 -56 189
rect -25 180 -23 182
rect -90 161 -88 163
rect -82 159 -80 163
rect -74 161 -72 163
rect -103 157 -80 159
rect -77 159 -72 161
rect -103 140 -101 157
rect -85 149 -83 154
rect -77 149 -75 159
rect -66 158 -64 163
rect -58 161 -56 163
rect -25 162 -23 172
rect -38 161 -37 162
rect -69 157 -64 158
rect -73 156 -64 157
rect -62 159 -37 161
rect -73 155 -67 156
rect -73 149 -71 155
rect -62 154 -60 159
rect -38 158 -37 159
rect -33 158 -23 162
rect -25 156 -23 158
rect 55 163 57 221
rect 55 161 158 163
rect -65 152 -60 154
rect -65 149 -63 152
rect -58 149 -56 151
rect -25 150 -23 152
rect 55 149 57 161
rect 80 157 82 161
rect 156 159 183 161
rect 88 157 90 159
rect 96 157 98 159
rect -129 138 -101 140
rect -129 136 -127 138
rect 156 149 158 159
rect 181 157 183 159
rect 189 157 191 159
rect 197 157 199 159
rect -85 135 -83 137
rect -129 112 -127 128
rect -77 114 -75 137
rect -73 135 -71 137
rect -65 135 -63 137
rect -58 135 -56 137
rect -61 133 -56 135
rect -129 106 -127 108
rect -61 106 -59 133
rect 55 125 57 141
rect 80 139 82 141
rect 88 130 90 141
rect 83 126 85 130
rect 88 128 92 130
rect 83 124 88 126
rect 86 122 88 124
rect 90 122 92 128
rect 96 125 98 141
rect 156 125 158 141
rect 181 139 183 141
rect 189 130 191 141
rect 185 126 187 130
rect 189 128 193 130
rect 94 123 98 125
rect 94 122 96 123
rect 55 119 57 121
rect 185 124 189 126
rect 187 122 189 124
rect 191 122 193 128
rect 197 125 199 141
rect 195 123 199 125
rect 195 122 197 123
rect 86 108 88 110
rect -129 104 39 106
rect 12 102 14 104
rect 37 96 39 104
rect 90 96 92 110
rect 37 94 92 96
rect 12 84 14 90
rect 94 87 96 110
rect 94 85 101 87
rect -142 80 14 84
rect 12 78 14 80
rect -56 69 -54 72
rect -142 65 -54 69
rect -64 44 -62 46
rect -56 44 -54 65
rect -48 44 -46 72
rect 12 70 14 72
rect 83 65 85 67
rect 91 65 93 67
rect 99 65 101 85
rect 156 69 158 121
rect 187 108 189 110
rect 191 92 193 110
rect 195 92 197 110
rect 156 67 183 69
rect 58 57 60 59
rect 156 57 158 67
rect 181 65 183 67
rect 189 65 191 67
rect 197 65 199 67
rect 58 47 60 49
rect 83 47 85 49
rect 58 45 85 47
rect -91 36 -89 38
rect -18 36 -16 38
rect 58 33 60 45
rect 91 38 93 49
rect 87 34 89 38
rect 91 36 95 38
rect 87 32 91 34
rect 89 30 91 32
rect 93 30 95 36
rect 99 33 101 49
rect 156 33 158 49
rect 181 47 183 49
rect 189 38 191 49
rect 185 34 187 38
rect 189 36 193 38
rect 97 31 101 33
rect 97 30 99 31
rect -91 26 -89 28
rect -64 26 -62 28
rect -91 24 -62 26
rect -91 19 -89 24
rect -97 15 -89 19
rect -56 17 -54 28
rect -91 12 -89 15
rect -65 13 -63 17
rect -56 15 -52 17
rect -65 11 -56 13
rect -58 9 -56 11
rect -54 9 -52 15
rect -48 12 -46 28
rect -18 18 -16 28
rect -26 14 -16 18
rect -18 12 -16 14
rect -50 10 -46 12
rect -50 9 -48 10
rect -91 -16 -89 8
rect -18 6 -16 8
rect -58 -5 -56 -3
rect -54 -5 -52 -3
rect -50 -5 -48 -3
rect 58 -16 60 29
rect 185 32 189 34
rect 187 30 189 32
rect 191 30 193 36
rect 197 33 199 49
rect 195 31 199 33
rect 195 30 197 31
rect 89 16 91 18
rect 93 0 95 18
rect 97 -7 99 18
rect 156 -16 158 29
rect 187 16 189 18
rect 191 0 193 18
rect 195 0 197 18
rect -91 -18 158 -16
<< ndiffusion >>
rect -141 191 -139 195
rect -135 191 -134 195
rect -132 191 -131 195
rect -127 191 -125 195
rect -32 152 -30 156
rect -26 152 -25 156
rect -23 152 -22 156
rect -18 152 -16 156
rect -95 143 -85 149
rect -95 139 -90 143
rect -86 139 -85 143
rect -95 137 -85 139
rect -83 142 -77 149
rect -83 138 -82 142
rect -78 138 -77 142
rect -83 137 -77 138
rect -75 137 -73 149
rect -71 145 -70 149
rect -66 145 -65 149
rect -71 137 -65 145
rect -63 137 -58 149
rect -56 142 -51 149
rect -56 138 -55 142
rect -56 137 -51 138
rect -136 108 -134 112
rect -130 108 -129 112
rect -127 108 -126 112
rect -122 108 -120 112
rect 49 121 50 125
rect 54 121 55 125
rect 57 121 58 125
rect 62 121 63 125
rect 80 116 86 122
rect 80 112 81 116
rect 85 112 86 116
rect 80 110 86 112
rect 88 110 90 122
rect 92 110 94 122
rect 96 116 103 122
rect 150 121 151 125
rect 155 121 156 125
rect 158 121 159 125
rect 163 121 164 125
rect 96 112 97 116
rect 101 112 103 116
rect 96 110 103 112
rect 5 74 7 78
rect 11 74 12 78
rect 5 72 12 74
rect 14 74 15 78
rect 19 74 21 78
rect 14 72 21 74
rect 181 116 187 122
rect 181 112 182 116
rect 186 112 187 116
rect 181 110 187 112
rect 189 110 191 122
rect 193 110 195 122
rect 197 116 204 122
rect 197 112 198 116
rect 202 112 204 116
rect 197 110 204 112
rect 52 29 53 33
rect 57 29 58 33
rect 60 29 61 33
rect 65 29 66 33
rect -97 8 -96 12
rect -92 8 -91 12
rect -89 8 -88 12
rect -84 8 -83 12
rect -64 3 -58 9
rect -64 -1 -63 3
rect -59 -1 -58 3
rect -64 -3 -58 -1
rect -56 -3 -54 9
rect -52 -3 -50 9
rect -48 3 -41 9
rect -24 8 -23 12
rect -19 8 -18 12
rect -16 8 -15 12
rect -11 8 -10 12
rect -48 -1 -47 3
rect -43 -1 -41 3
rect -48 -3 -41 -1
rect 83 24 89 30
rect 83 20 84 24
rect 88 20 89 24
rect 83 18 89 20
rect 91 18 93 30
rect 95 18 97 30
rect 99 24 106 30
rect 150 29 151 33
rect 155 29 156 33
rect 158 29 159 33
rect 163 29 164 33
rect 99 20 100 24
rect 104 20 106 24
rect 99 18 106 20
rect 181 24 187 30
rect 181 20 182 24
rect 186 20 187 24
rect 181 18 187 20
rect 189 18 191 30
rect 193 18 195 30
rect 197 24 204 30
rect 197 20 198 24
rect 202 20 204 24
rect 197 18 204 20
<< pdiffusion >>
rect -140 215 -139 219
rect -135 215 -134 219
rect -140 211 -134 215
rect -132 215 -131 219
rect -127 215 -126 219
rect -132 211 -126 215
rect -95 183 -90 187
rect -91 179 -90 183
rect -95 163 -90 179
rect -88 182 -82 187
rect -88 178 -87 182
rect -83 178 -82 182
rect -88 163 -82 178
rect -80 175 -74 187
rect -80 171 -79 175
rect -75 171 -74 175
rect -80 163 -74 171
rect -72 167 -66 187
rect -72 163 -71 167
rect -67 163 -66 167
rect -64 175 -58 187
rect -64 171 -63 175
rect -59 171 -58 175
rect -64 163 -58 171
rect -56 182 -51 187
rect -56 178 -55 182
rect -56 163 -51 178
rect -31 176 -30 180
rect -26 176 -25 180
rect -31 172 -25 176
rect -23 176 -22 180
rect -18 176 -17 180
rect -23 172 -17 176
rect 75 156 80 157
rect 79 152 80 156
rect 49 145 50 149
rect 54 145 55 149
rect 49 141 55 145
rect 57 145 58 149
rect 62 145 63 149
rect 57 141 63 145
rect 75 141 80 152
rect 82 156 88 157
rect 82 152 83 156
rect 87 152 88 156
rect 82 141 88 152
rect 90 147 96 157
rect 90 143 91 147
rect 95 143 96 147
rect 90 141 96 143
rect 98 156 103 157
rect 98 152 99 156
rect 98 141 103 152
rect 176 156 181 157
rect 180 152 181 156
rect 150 145 151 149
rect 155 145 156 149
rect 150 141 156 145
rect 158 145 159 149
rect 163 145 164 149
rect 158 141 164 145
rect 176 141 181 152
rect 183 156 189 157
rect 183 152 184 156
rect 188 152 189 156
rect 183 141 189 152
rect 191 147 197 157
rect 191 143 192 147
rect 196 143 197 147
rect 191 141 197 143
rect 199 156 204 157
rect 199 152 200 156
rect 199 141 204 152
rect -135 132 -134 136
rect -130 132 -129 136
rect -135 128 -129 132
rect -127 132 -126 136
rect -122 132 -121 136
rect -127 128 -121 132
rect 6 98 7 102
rect 11 98 12 102
rect 6 90 12 98
rect 14 98 15 102
rect 19 98 20 102
rect 14 90 20 98
rect 78 64 83 65
rect 82 60 83 64
rect 52 53 53 57
rect 57 53 58 57
rect 52 49 58 53
rect 60 53 61 57
rect 65 53 66 57
rect 60 49 66 53
rect 78 49 83 60
rect 85 64 91 65
rect 85 60 86 64
rect 90 60 91 64
rect 85 49 91 60
rect 93 55 99 65
rect 93 51 94 55
rect 98 51 99 55
rect 93 49 99 51
rect 101 64 106 65
rect 101 60 102 64
rect 101 49 106 60
rect 176 64 181 65
rect 180 60 181 64
rect 150 53 151 57
rect 155 53 156 57
rect 150 49 156 53
rect 158 53 159 57
rect 163 53 164 57
rect 158 49 164 53
rect 176 49 181 60
rect 183 64 189 65
rect 183 60 184 64
rect 188 60 189 64
rect 183 49 189 60
rect 191 55 197 65
rect 191 51 192 55
rect 196 51 197 55
rect 191 49 197 51
rect 199 64 204 65
rect 199 60 200 64
rect 199 49 204 60
rect -69 43 -64 44
rect -65 39 -64 43
rect -97 32 -96 36
rect -92 32 -91 36
rect -97 28 -91 32
rect -89 32 -88 36
rect -84 32 -83 36
rect -89 28 -83 32
rect -69 28 -64 39
rect -62 43 -56 44
rect -62 39 -61 43
rect -57 39 -56 43
rect -62 28 -56 39
rect -54 34 -48 44
rect -54 30 -53 34
rect -49 30 -48 34
rect -54 28 -48 30
rect -46 43 -41 44
rect -46 39 -45 43
rect -46 28 -41 39
rect -24 32 -23 36
rect -19 32 -18 36
rect -24 28 -18 32
rect -16 32 -15 36
rect -11 32 -10 36
rect -16 28 -10 32
<< metal1 >>
rect -143 239 -123 241
rect -143 235 -139 239
rect -135 235 -123 239
rect -143 233 -123 235
rect -139 219 -135 233
rect -131 201 -127 215
rect -41 207 -3 211
rect -131 197 -105 201
rect -131 195 -127 197
rect -139 177 -135 191
rect -143 176 -123 177
rect -143 172 -139 176
rect -135 172 -123 176
rect -143 169 -123 172
rect -138 156 -118 158
rect -138 152 -134 156
rect -130 152 -118 156
rect -138 150 -118 152
rect -109 154 -105 197
rect -99 199 -55 201
rect -99 195 -95 199
rect -91 195 -55 199
rect -99 193 -55 195
rect -34 200 -14 202
rect -34 196 -30 200
rect -26 196 -14 200
rect -34 194 -14 196
rect -95 183 -91 193
rect -83 178 -55 182
rect -30 180 -26 194
rect -75 171 -63 175
rect -71 158 -67 163
rect -22 162 -18 176
rect -7 162 -3 207
rect -71 155 -44 158
rect -70 154 -44 155
rect -109 150 -89 154
rect -134 136 -130 150
rect -70 149 -66 154
rect -90 132 -86 139
rect -78 138 -55 142
rect -126 118 -122 132
rect -100 130 -56 132
rect -100 126 -90 130
rect -86 126 -56 130
rect -100 124 -56 126
rect -126 114 -81 118
rect -126 112 -122 114
rect -134 94 -130 108
rect -48 103 -44 154
rect -37 144 -33 158
rect -22 158 -3 162
rect 19 174 230 178
rect -22 156 -18 158
rect -41 141 -33 144
rect -41 126 -37 141
rect -30 138 -26 152
rect -34 137 -14 138
rect -34 133 -30 137
rect -26 133 -14 137
rect 19 136 23 174
rect 46 169 112 171
rect 46 165 50 169
rect 54 165 75 169
rect 79 165 99 169
rect 103 165 112 169
rect 46 163 112 165
rect 147 169 213 171
rect 147 165 151 169
rect 155 165 176 169
rect 180 165 200 169
rect 204 165 213 169
rect 147 163 213 165
rect 50 149 54 163
rect 75 156 79 163
rect 87 152 99 156
rect 151 149 155 163
rect 176 156 180 163
rect 188 152 200 156
rect -34 130 -14 133
rect -8 132 23 136
rect -8 126 -4 132
rect -41 122 -4 126
rect 58 130 62 145
rect 91 138 95 143
rect 91 134 109 138
rect 105 131 109 134
rect 58 126 79 130
rect 105 127 135 131
rect 58 125 62 126
rect 3 122 23 124
rect 3 118 7 122
rect 11 118 23 122
rect 3 116 23 118
rect -48 99 -42 103
rect -138 93 -118 94
rect -138 89 -134 93
rect -130 89 -118 93
rect -138 86 -118 89
rect -46 69 -42 99
rect 7 102 11 116
rect 50 107 54 121
rect 105 116 109 127
rect 101 112 109 116
rect 81 107 85 112
rect 46 106 112 107
rect 46 102 50 106
rect 54 105 112 106
rect 54 102 81 105
rect 46 101 81 102
rect 85 101 112 105
rect 46 99 112 101
rect 15 84 19 98
rect 131 96 135 127
rect 159 130 163 145
rect 192 138 196 143
rect 192 134 210 138
rect 206 130 210 134
rect 226 130 230 174
rect 159 126 181 130
rect 206 126 234 130
rect 159 125 163 126
rect 151 107 155 121
rect 206 116 210 126
rect 202 112 210 116
rect 182 107 186 112
rect 147 106 213 107
rect 147 102 151 106
rect 155 105 213 106
rect 155 102 182 105
rect 147 101 182 102
rect 186 101 213 105
rect 147 99 213 101
rect 131 92 187 96
rect 201 92 220 96
rect 15 80 38 84
rect 15 78 19 80
rect 7 60 11 74
rect 3 59 23 60
rect -100 56 -7 58
rect -100 52 -96 56
rect -92 52 -69 56
rect -65 52 -45 56
rect -41 52 -23 56
rect -19 52 -7 56
rect 3 55 7 59
rect 11 55 23 59
rect 3 52 23 55
rect -100 50 -7 52
rect -96 36 -92 50
rect -69 43 -65 50
rect -57 39 -45 43
rect -23 36 -19 50
rect -88 17 -84 32
rect -53 25 -49 30
rect -53 21 -35 25
rect -39 18 -35 21
rect -15 18 -11 32
rect -88 13 -69 17
rect -39 14 -30 18
rect -39 13 -26 14
rect -15 14 10 18
rect -88 12 -84 13
rect -96 -6 -92 8
rect -39 3 -35 13
rect -15 12 -11 14
rect -43 -1 -35 3
rect -63 -6 -59 -1
rect -23 -6 -19 8
rect 6 -3 10 14
rect 34 4 38 80
rect 49 77 115 79
rect 49 73 53 77
rect 57 73 78 77
rect 82 73 102 77
rect 106 73 115 77
rect 49 71 115 73
rect 147 77 213 79
rect 147 73 151 77
rect 155 73 176 77
rect 180 73 200 77
rect 204 73 213 77
rect 147 71 213 73
rect 53 57 57 71
rect 78 64 82 71
rect 90 60 102 64
rect 151 57 155 71
rect 176 64 180 71
rect 188 60 200 64
rect 61 38 65 53
rect 94 46 98 51
rect 94 42 112 46
rect 108 39 112 42
rect 61 34 83 38
rect 108 35 133 39
rect 61 33 65 34
rect 53 15 57 29
rect 108 24 112 35
rect 104 20 112 24
rect 84 15 88 20
rect 49 14 115 15
rect 49 10 53 14
rect 57 13 115 14
rect 57 10 84 13
rect 49 9 84 10
rect 88 9 115 13
rect 49 7 115 9
rect 129 4 133 35
rect 159 38 163 53
rect 192 46 196 51
rect 192 42 210 46
rect 206 39 210 42
rect 216 39 220 92
rect 159 34 181 38
rect 206 35 220 39
rect 159 33 163 34
rect 151 15 155 29
rect 206 24 210 35
rect 202 20 210 24
rect 182 15 186 20
rect 147 14 213 15
rect 147 10 151 14
rect 155 13 213 14
rect 155 10 182 13
rect 147 9 182 10
rect 186 9 213 13
rect 147 7 213 9
rect 226 4 230 126
rect 34 0 89 4
rect 129 0 187 4
rect 201 0 230 4
rect -100 -7 -7 -6
rect 6 -7 93 -3
rect -100 -11 -96 -7
rect -92 -8 -23 -7
rect -92 -11 -63 -8
rect -100 -12 -63 -11
rect -59 -11 -23 -8
rect -19 -11 -7 -7
rect -59 -12 -7 -11
rect -100 -14 -7 -12
<< ntransistor >>
rect -134 191 -132 195
rect -25 152 -23 156
rect -85 137 -83 149
rect -77 137 -75 149
rect -73 137 -71 149
rect -65 137 -63 149
rect -58 137 -56 149
rect -129 108 -127 112
rect 55 121 57 125
rect 86 110 88 122
rect 90 110 92 122
rect 94 110 96 122
rect 156 121 158 125
rect 12 72 14 78
rect 187 110 189 122
rect 191 110 193 122
rect 195 110 197 122
rect 58 29 60 33
rect -91 8 -89 12
rect -58 -3 -56 9
rect -54 -3 -52 9
rect -50 -3 -48 9
rect -18 8 -16 12
rect 89 18 91 30
rect 93 18 95 30
rect 97 18 99 30
rect 156 29 158 33
rect 187 18 189 30
rect 191 18 193 30
rect 195 18 197 30
<< ptransistor >>
rect -134 211 -132 219
rect -90 163 -88 187
rect -82 163 -80 187
rect -74 163 -72 187
rect -66 163 -64 187
rect -58 163 -56 187
rect -25 172 -23 180
rect 55 141 57 149
rect 80 141 82 157
rect 88 141 90 157
rect 96 141 98 157
rect 156 141 158 149
rect 181 141 183 157
rect 189 141 191 157
rect 197 141 199 157
rect -129 128 -127 136
rect 12 90 14 102
rect 58 49 60 57
rect 83 49 85 65
rect 91 49 93 65
rect 99 49 101 65
rect 156 49 158 57
rect 181 49 183 65
rect 189 49 191 65
rect 197 49 199 65
rect -91 28 -89 36
rect -64 28 -62 44
rect -56 28 -54 44
rect -48 28 -46 44
rect -18 28 -16 36
<< polycontact >>
rect -146 197 -142 201
rect -45 207 -41 211
rect -89 150 -85 154
rect -37 158 -33 162
rect -81 114 -77 118
rect 79 126 83 130
rect 181 126 185 130
rect -146 80 -142 84
rect -146 65 -142 69
rect -46 65 -42 69
rect 187 92 191 96
rect 197 92 201 96
rect 83 34 87 38
rect 181 34 185 38
rect -101 15 -97 19
rect -69 13 -65 17
rect -30 14 -26 18
rect 89 0 93 4
rect 93 -7 97 -3
rect 187 0 191 4
rect 197 0 201 4
<< ndcontact >>
rect -139 191 -135 195
rect -131 191 -127 195
rect -30 152 -26 156
rect -22 152 -18 156
rect -90 139 -86 143
rect -82 138 -78 142
rect -70 145 -66 149
rect -55 138 -51 142
rect -134 108 -130 112
rect -126 108 -122 112
rect 50 121 54 125
rect 58 121 62 125
rect 81 112 85 116
rect 151 121 155 125
rect 159 121 163 125
rect 97 112 101 116
rect 7 74 11 78
rect 15 74 19 78
rect 182 112 186 116
rect 198 112 202 116
rect 53 29 57 33
rect 61 29 65 33
rect -96 8 -92 12
rect -88 8 -84 12
rect -63 -1 -59 3
rect -23 8 -19 12
rect -15 8 -11 12
rect -47 -1 -43 3
rect 84 20 88 24
rect 151 29 155 33
rect 159 29 163 33
rect 100 20 104 24
rect 182 20 186 24
rect 198 20 202 24
<< pdcontact >>
rect -139 215 -135 219
rect -131 215 -127 219
rect -95 179 -91 183
rect -87 178 -83 182
rect -79 171 -75 175
rect -71 163 -67 167
rect -63 171 -59 175
rect -55 178 -51 182
rect -30 176 -26 180
rect -22 176 -18 180
rect 75 152 79 156
rect 50 145 54 149
rect 58 145 62 149
rect 83 152 87 156
rect 91 143 95 147
rect 99 152 103 156
rect 176 152 180 156
rect 151 145 155 149
rect 159 145 163 149
rect 184 152 188 156
rect 192 143 196 147
rect 200 152 204 156
rect -134 132 -130 136
rect -126 132 -122 136
rect 7 98 11 102
rect 15 98 19 102
rect 78 60 82 64
rect 53 53 57 57
rect 61 53 65 57
rect 86 60 90 64
rect 94 51 98 55
rect 102 60 106 64
rect 176 60 180 64
rect 151 53 155 57
rect 159 53 163 57
rect 184 60 188 64
rect 192 51 196 55
rect 200 60 204 64
rect -69 39 -65 43
rect -96 32 -92 36
rect -88 32 -84 36
rect -61 39 -57 43
rect -53 30 -49 34
rect -45 39 -41 43
rect -23 32 -19 36
rect -15 32 -11 36
<< psubstratepcontact >>
rect -139 172 -135 176
rect -90 126 -86 130
rect -30 133 -26 137
rect -134 89 -130 93
rect 50 102 54 106
rect 81 101 85 105
rect 151 102 155 106
rect 182 101 186 105
rect 7 55 11 59
rect -96 -11 -92 -7
rect 53 10 57 14
rect -63 -12 -59 -8
rect -23 -11 -19 -7
rect 84 9 88 13
rect 151 10 155 14
rect 182 9 186 13
<< nsubstratencontact >>
rect -139 235 -135 239
rect -95 195 -91 199
rect -30 196 -26 200
rect -134 152 -130 156
rect 50 165 54 169
rect 75 165 79 169
rect 99 165 103 169
rect 151 165 155 169
rect 176 165 180 169
rect 200 165 204 169
rect 7 118 11 122
rect 53 73 57 77
rect 78 73 82 77
rect -96 52 -92 56
rect -69 52 -65 56
rect 102 73 106 77
rect 151 73 155 77
rect 176 73 180 77
rect 200 73 204 77
rect -45 52 -41 56
rect -23 52 -19 56
<< labels >>
rlabel metal1 19 80 22 84 5 d_n
rlabel nwell 46 163 112 171 1 vdd_1
rlabel nwell 147 163 213 171 1 vdd_2
rlabel nwell 147 71 213 79 1 vdd_4
rlabel nwell 49 71 115 79 1 vdd_3
rlabel metal1 46 99 112 107 5 vss_1
rlabel metal1 147 99 213 107 5 vss_2
rlabel metal1 147 7 213 15 5 vss_4
rlabel metal1 49 7 115 15 5 vss_3
rlabel metal1 230 126 234 130 3 out
rlabel polycontact 93 -7 97 -3 5 gated_clk
rlabel metal1 3 52 23 60 5 vss_5
rlabel nwell 3 116 23 124 1 vdd_5
rlabel nwell -100 50 -7 58 1 vdd_10
rlabel metal1 -100 -14 -7 -6 5 vss_10
rlabel polycontact -101 15 -97 19 7 sleep
rlabel polycontact -146 197 -142 201 5 sleep
rlabel nwell -143 233 -123 241 1 vdd_6
rlabel metal1 -143 169 -123 177 5 vss_6
rlabel nwell -138 150 -118 158 1 vdd_7
rlabel metal1 -138 86 -118 94 5 vss_7
rlabel metal1 -99 193 -55 201 1 vdd_8
rlabel metal1 -100 124 -56 132 5 vss_8
rlabel nwell -34 194 -14 202 1 vdd_9
rlabel metal1 -34 130 -14 138 5 vss_9
rlabel polycontact -146 80 -142 84 7 d
rlabel polycontact -146 65 -142 69 7 clk
<< end >>
