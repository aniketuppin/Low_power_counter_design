magic
tech scmos
timestamp 1678956533
<< nwell >>
rect -11 111 16 149
rect 34 70 90 107
rect 99 72 125 113
rect -6 28 21 69
<< polysilicon >>
rect 1 127 3 129
rect 88 119 94 120
rect 1 109 3 119
rect -7 105 3 109
rect 88 115 90 119
rect 88 114 94 115
rect 1 103 3 105
rect 88 101 90 114
rect 69 99 90 101
rect 1 97 3 99
rect 23 97 47 99
rect 1 95 25 97
rect 45 95 47 97
rect 53 95 55 97
rect 61 95 63 97
rect 69 95 71 99
rect 77 95 79 97
rect 110 88 112 90
rect 45 69 47 71
rect 53 67 55 71
rect 61 69 63 71
rect 32 65 55 67
rect 58 67 63 69
rect 32 48 34 65
rect 50 57 52 62
rect 58 57 60 67
rect 69 66 71 71
rect 77 69 79 71
rect 110 70 112 80
rect 97 69 98 70
rect 66 65 71 66
rect 62 64 71 65
rect 73 67 98 69
rect 62 63 68 64
rect 62 57 64 63
rect 73 62 75 67
rect 97 66 98 67
rect 102 66 112 70
rect 110 64 112 66
rect 70 60 75 62
rect 70 57 72 60
rect 77 57 79 59
rect 110 58 112 60
rect 6 46 34 48
rect 6 44 8 46
rect 50 43 52 45
rect 6 26 8 36
rect -2 22 8 26
rect 58 22 60 45
rect 62 43 64 45
rect 70 43 72 45
rect 77 43 79 45
rect 74 41 79 43
rect 6 20 8 22
rect 6 14 8 16
rect 74 14 76 41
rect 6 12 76 14
<< ndiffusion >>
rect -6 99 -4 103
rect 0 99 1 103
rect 3 99 4 103
rect 8 99 10 103
rect 103 60 105 64
rect 109 60 110 64
rect 112 60 113 64
rect 117 60 119 64
rect 40 51 50 57
rect 40 47 45 51
rect 49 47 50 51
rect 40 45 50 47
rect 52 50 58 57
rect 52 46 53 50
rect 57 46 58 50
rect 52 45 58 46
rect 60 45 62 57
rect 64 53 65 57
rect 69 53 70 57
rect 64 45 70 53
rect 72 45 77 57
rect 79 50 84 57
rect 79 46 80 50
rect 79 45 84 46
rect -1 16 1 20
rect 5 16 6 20
rect 8 16 9 20
rect 13 16 15 20
<< pdiffusion >>
rect -5 123 -4 127
rect 0 123 1 127
rect -5 119 1 123
rect 3 123 4 127
rect 8 123 9 127
rect 3 119 9 123
rect 40 91 45 95
rect 44 87 45 91
rect 40 71 45 87
rect 47 90 53 95
rect 47 86 48 90
rect 52 86 53 90
rect 47 71 53 86
rect 55 83 61 95
rect 55 79 56 83
rect 60 79 61 83
rect 55 71 61 79
rect 63 75 69 95
rect 63 71 64 75
rect 68 71 69 75
rect 71 83 77 95
rect 71 79 72 83
rect 76 79 77 83
rect 71 71 77 79
rect 79 90 84 95
rect 79 86 80 90
rect 79 71 84 86
rect 104 84 105 88
rect 109 84 110 88
rect 104 80 110 84
rect 112 84 113 88
rect 117 84 118 88
rect 112 80 118 84
rect 0 40 1 44
rect 5 40 6 44
rect 0 36 6 40
rect 8 40 9 44
rect 13 40 14 44
rect 8 36 14 40
<< metal1 >>
rect -8 147 12 149
rect -8 143 -4 147
rect 0 143 12 147
rect -8 141 12 143
rect -4 127 0 141
rect 4 109 8 123
rect 94 115 132 119
rect 4 105 30 109
rect 4 103 8 105
rect -4 85 0 99
rect -8 84 12 85
rect -8 80 -4 84
rect 0 80 12 84
rect -8 77 12 80
rect -3 64 17 66
rect -3 60 1 64
rect 5 60 17 64
rect -3 58 17 60
rect 26 62 30 105
rect 36 107 80 109
rect 36 103 40 107
rect 44 103 80 107
rect 36 101 80 103
rect 101 108 121 110
rect 101 104 105 108
rect 109 104 121 108
rect 101 102 121 104
rect 40 91 44 101
rect 52 86 80 90
rect 105 88 109 102
rect 60 79 72 83
rect 64 66 68 71
rect 113 70 117 84
rect 128 70 132 115
rect 113 66 132 70
rect 64 63 89 66
rect 113 64 117 66
rect 65 62 89 63
rect 26 58 46 62
rect 1 44 5 58
rect 65 57 69 62
rect 45 40 49 47
rect 57 46 80 50
rect 105 46 109 60
rect 101 45 121 46
rect 101 41 105 45
rect 109 41 121 45
rect 9 26 13 40
rect 35 38 79 40
rect 101 38 121 41
rect 35 34 45 38
rect 49 34 79 38
rect 35 32 79 34
rect 9 22 54 26
rect 9 20 13 22
rect 1 2 5 16
rect -3 1 17 2
rect -3 -3 1 1
rect 5 -3 17 1
rect -3 -6 17 -3
<< ntransistor >>
rect 1 99 3 103
rect 110 60 112 64
rect 50 45 52 57
rect 58 45 60 57
rect 62 45 64 57
rect 70 45 72 57
rect 77 45 79 57
rect 6 16 8 20
<< ptransistor >>
rect 1 119 3 127
rect 45 71 47 95
rect 53 71 55 95
rect 61 71 63 95
rect 69 71 71 95
rect 77 71 79 95
rect 110 80 112 88
rect 6 36 8 44
<< polycontact >>
rect -11 105 -7 109
rect 90 115 94 119
rect 46 58 50 62
rect 98 66 102 70
rect -6 22 -2 26
rect 54 22 58 26
<< ndcontact >>
rect -4 99 0 103
rect 4 99 8 103
rect 105 60 109 64
rect 113 60 117 64
rect 45 47 49 51
rect 53 46 57 50
rect 65 53 69 57
rect 80 46 84 50
rect 1 16 5 20
rect 9 16 13 20
<< pdcontact >>
rect -4 123 0 127
rect 4 123 8 127
rect 40 87 44 91
rect 48 86 52 90
rect 56 79 60 83
rect 64 71 68 75
rect 72 79 76 83
rect 80 86 84 90
rect 105 84 109 88
rect 113 84 117 88
rect 1 40 5 44
rect 9 40 13 44
<< psubstratepcontact >>
rect -4 80 0 84
rect 45 34 49 38
rect 105 41 109 45
rect 1 -3 5 1
<< nsubstratencontact >>
rect -4 143 0 147
rect 40 103 44 107
rect 105 104 109 108
rect 1 60 5 64
<< labels >>
rlabel polycontact 98 66 102 70 5 a
rlabel polycontact -6 22 -2 26 5 b
rlabel metal1 85 62 89 66 3 out
rlabel metal1 35 32 79 40 1 vss
rlabel polycontact -11 105 -7 109 5 sleep
rlabel metal1 36 101 80 109 1 vdd
rlabel metal1 101 38 121 46 1 vss_3
rlabel metal1 -3 -6 17 2 5 vss_2
rlabel nwell -3 58 17 66 1 vdd_2
rlabel metal1 -8 77 12 85 5 vss_1
rlabel nwell -8 141 12 149 1 vdd_1
rlabel nwell 101 102 121 110 1 vdd_3
<< end >>
