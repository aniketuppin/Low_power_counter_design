magic
tech scmos
timestamp 1678735475
<< nwell >>
rect -39 72 -12 75
rect 34 72 61 75
rect -39 41 61 72
rect -39 34 -12 41
rect 34 34 61 41
<< polysilicon >>
rect 0 58 2 60
rect 8 58 10 60
rect 16 58 18 60
rect -27 50 -25 52
rect 46 50 48 52
rect -27 40 -25 42
rect 0 40 2 42
rect -27 38 2 40
rect -27 32 -25 38
rect -35 28 -25 32
rect 8 31 10 42
rect 16 32 18 42
rect 46 32 48 42
rect 16 31 23 32
rect -27 26 -25 28
rect -1 27 1 31
rect 8 29 12 31
rect -1 25 8 27
rect 6 23 8 25
rect 10 23 12 29
rect 16 27 18 31
rect 22 27 23 31
rect 38 28 48 32
rect 16 26 23 27
rect 46 26 48 28
rect 14 24 18 26
rect 14 23 16 24
rect -27 20 -25 22
rect 46 20 48 22
rect 6 9 8 11
rect 10 9 12 11
rect 14 9 16 11
<< ndiffusion >>
rect -33 22 -32 26
rect -28 22 -27 26
rect -25 22 -24 26
rect -20 22 -19 26
rect 0 17 6 23
rect 0 13 1 17
rect 5 13 6 17
rect 0 11 6 13
rect 8 11 10 23
rect 12 11 14 23
rect 16 17 23 23
rect 40 22 41 26
rect 45 22 46 26
rect 48 22 49 26
rect 53 22 54 26
rect 16 13 17 17
rect 21 13 23 17
rect 16 11 23 13
<< pdiffusion >>
rect -5 57 0 58
rect -1 53 0 57
rect -33 46 -32 50
rect -28 46 -27 50
rect -33 42 -27 46
rect -25 46 -24 50
rect -20 46 -19 50
rect -25 42 -19 46
rect -5 42 0 53
rect 2 57 8 58
rect 2 53 3 57
rect 7 53 8 57
rect 2 42 8 53
rect 10 48 16 58
rect 10 44 11 48
rect 15 44 16 48
rect 10 42 16 44
rect 18 57 23 58
rect 18 53 19 57
rect 18 42 23 53
rect 40 46 41 50
rect 45 46 46 50
rect 40 42 46 46
rect 48 46 49 50
rect 53 46 54 50
rect 48 42 54 46
<< metal1 >>
rect -36 70 57 72
rect -36 66 -32 70
rect -28 66 -5 70
rect -1 66 19 70
rect 23 66 41 70
rect 45 66 57 70
rect -36 64 57 66
rect -32 50 -28 64
rect -5 57 -1 64
rect 7 53 19 57
rect 41 50 45 64
rect -24 31 -20 46
rect 11 39 15 44
rect 11 35 29 39
rect 25 32 29 35
rect 49 32 53 46
rect -24 27 -5 31
rect 25 28 34 32
rect 25 27 38 28
rect 49 28 56 32
rect -24 26 -20 27
rect -32 8 -28 22
rect 25 17 29 27
rect 49 26 53 28
rect 21 13 29 17
rect 1 8 5 13
rect 41 8 45 22
rect -36 7 57 8
rect -36 3 -32 7
rect -28 6 41 7
rect -28 3 1 6
rect -36 2 1 3
rect 5 3 41 6
rect 45 3 57 7
rect 5 2 57 3
rect -36 0 57 2
<< ntransistor >>
rect -27 22 -25 26
rect 6 11 8 23
rect 10 11 12 23
rect 14 11 16 23
rect 46 22 48 26
<< ptransistor >>
rect -27 42 -25 50
rect 0 42 2 58
rect 8 42 10 58
rect 16 42 18 58
rect 46 42 48 50
<< polycontact >>
rect -39 28 -35 32
rect 4 31 8 35
rect -5 27 -1 31
rect 18 27 22 31
rect 34 28 38 32
<< ndcontact >>
rect -32 22 -28 26
rect -24 22 -20 26
rect 1 13 5 17
rect 41 22 45 26
rect 49 22 53 26
rect 17 13 21 17
<< pdcontact >>
rect -5 53 -1 57
rect -32 46 -28 50
rect -24 46 -20 50
rect 3 53 7 57
rect 11 44 15 48
rect 19 53 23 57
rect 41 46 45 50
rect 49 46 53 50
<< psubstratepcontact >>
rect -32 3 -28 7
rect 1 2 5 6
rect 41 3 45 7
<< nsubstratencontact >>
rect -32 66 -28 70
rect -5 66 -1 70
rect 19 66 23 70
rect 41 66 45 70
<< labels >>
rlabel polycontact 18 27 22 31 5 b
rlabel polycontact -39 28 -35 32 7 sleep
rlabel metal1 53 28 56 32 3 out
rlabel nwell -36 64 57 72 1 vdd
rlabel metal1 -36 0 57 8 5 vss
rlabel polycontact 4 31 8 35 5 a
<< end >>
