magic
tech scmos
timestamp 1679582807
<< nwell >>
rect -350 213 -281 244
rect -252 213 -183 244
rect -350 206 -323 213
rect -252 206 -225 213
rect -390 159 -363 200
rect -151 193 -124 231
rect 0 221 27 259
rect -106 152 -50 189
rect -41 154 -15 195
rect 45 180 101 217
rect 110 182 136 223
rect -350 121 -281 152
rect -252 121 -183 152
rect -350 114 -323 121
rect -252 114 -225 121
rect -146 110 -119 151
rect 5 138 32 179
rect 189 158 258 189
rect 290 158 359 189
rect 189 151 216 158
rect 290 151 317 158
rect 146 104 173 145
rect 43 76 70 79
rect 116 76 143 79
rect 43 45 143 76
rect 192 66 261 97
rect 290 66 359 97
rect 192 59 219 66
rect 290 59 317 66
rect 43 38 70 45
rect 116 38 143 45
<< polysilicon >>
rect -356 248 -197 250
rect -356 179 -354 248
rect -338 234 -238 236
rect -338 222 -336 234
rect -313 230 -311 234
rect -240 232 -213 234
rect -305 230 -303 232
rect -297 230 -295 232
rect -240 222 -238 232
rect -215 230 -213 232
rect -207 230 -205 232
rect -199 230 -197 248
rect -30 242 -26 243
rect -139 216 -66 218
rect -338 198 -336 214
rect -313 212 -311 214
rect -305 203 -303 214
rect -310 199 -308 203
rect -305 201 -301 203
rect -310 197 -305 199
rect -307 195 -305 197
rect -303 195 -301 201
rect -297 198 -295 214
rect -240 198 -238 214
rect -215 212 -213 214
rect -207 203 -205 214
rect -211 199 -209 203
rect -207 201 -203 203
rect -299 196 -295 198
rect -299 195 -297 196
rect -338 192 -336 194
rect -211 197 -207 199
rect -209 195 -207 197
rect -205 195 -203 201
rect -199 198 -197 214
rect -139 209 -137 216
rect -52 201 -46 202
rect -201 196 -197 198
rect -201 195 -199 196
rect -307 181 -305 183
rect -378 177 -354 179
rect -378 175 -376 177
rect -356 169 -354 177
rect -303 169 -301 183
rect -356 167 -301 169
rect -378 158 -376 163
rect -299 160 -297 183
rect -240 160 -238 194
rect -139 189 -137 201
rect -52 197 -50 201
rect -52 196 -46 197
rect -158 187 -137 189
rect -209 181 -207 183
rect -205 165 -203 183
rect -201 165 -199 183
rect -158 160 -156 187
rect -139 185 -137 187
rect -52 183 -50 196
rect -71 181 -50 183
rect -139 179 -137 181
rect -117 179 -93 181
rect -139 177 -115 179
rect -95 177 -93 179
rect -87 177 -85 179
rect -79 177 -77 179
rect -71 177 -69 181
rect -63 177 -61 179
rect -299 158 -295 160
rect -379 154 -376 158
rect -378 151 -376 154
rect -378 142 -376 145
rect -313 138 -311 140
rect -305 138 -303 140
rect -297 138 -295 158
rect -240 158 -156 160
rect -240 142 -238 158
rect -30 170 -28 242
rect 12 239 203 241
rect 12 237 14 239
rect 99 229 105 230
rect 12 219 14 229
rect 4 215 14 219
rect 99 225 101 229
rect 99 224 105 225
rect 12 213 14 215
rect 99 211 101 224
rect 80 209 101 211
rect 12 207 14 209
rect 34 207 58 209
rect 12 205 36 207
rect 56 205 58 207
rect 64 205 66 207
rect 72 205 74 207
rect 80 205 82 209
rect 88 205 90 207
rect 121 198 123 200
rect 56 179 58 181
rect 64 177 66 181
rect 72 179 74 181
rect 43 175 66 177
rect 69 177 74 179
rect -95 151 -93 153
rect -87 149 -85 153
rect -79 151 -77 153
rect -108 147 -85 149
rect -82 149 -77 151
rect -240 140 -213 142
rect -338 130 -336 132
rect -240 130 -238 140
rect -215 138 -213 140
rect -207 138 -205 140
rect -199 138 -197 140
rect -108 130 -106 147
rect -90 139 -88 144
rect -82 139 -80 149
rect -71 148 -69 153
rect -63 151 -61 153
rect -30 152 -28 162
rect 43 158 45 175
rect 61 167 63 172
rect 69 167 71 177
rect 80 176 82 181
rect 88 179 90 181
rect 121 180 123 190
rect 108 179 109 180
rect 77 175 82 176
rect 73 174 82 175
rect 84 177 109 179
rect 73 173 79 174
rect 73 167 75 173
rect 84 172 86 177
rect 108 176 109 177
rect 113 176 123 180
rect 121 174 123 176
rect 201 181 203 239
rect 201 179 304 181
rect 81 170 86 172
rect 81 167 83 170
rect 88 167 90 169
rect 121 168 123 170
rect 201 167 203 179
rect 226 175 228 179
rect 302 177 329 179
rect 234 175 236 177
rect 242 175 244 177
rect 17 156 45 158
rect 17 154 19 156
rect 302 167 304 177
rect 327 175 329 177
rect 335 175 337 177
rect 343 175 345 177
rect -43 151 -42 152
rect -74 147 -69 148
rect -78 146 -69 147
rect -67 149 -42 151
rect -78 145 -72 146
rect -78 139 -76 145
rect -67 144 -65 149
rect -43 148 -42 149
rect -38 148 -28 152
rect -30 146 -28 148
rect 61 153 63 155
rect -70 142 -65 144
rect -70 139 -68 142
rect -63 139 -61 141
rect -30 140 -28 142
rect -134 128 -106 130
rect -134 126 -132 128
rect 17 130 19 146
rect 69 132 71 155
rect 73 153 75 155
rect 81 153 83 155
rect 88 153 90 155
rect 85 151 90 153
rect -338 120 -336 122
rect -313 120 -311 122
rect -338 118 -311 120
rect -338 106 -336 118
rect -305 111 -303 122
rect -309 107 -307 111
rect -305 109 -301 111
rect -309 105 -305 107
rect -307 103 -305 105
rect -303 103 -301 109
rect -297 106 -295 122
rect -240 106 -238 122
rect -215 120 -213 122
rect -207 111 -205 122
rect -211 107 -209 111
rect -207 109 -203 111
rect -299 104 -295 106
rect -299 103 -297 104
rect -338 70 -336 102
rect -211 105 -207 107
rect -209 103 -207 105
rect -205 103 -203 109
rect -199 106 -197 122
rect -90 125 -88 127
rect -134 108 -132 118
rect -201 104 -197 106
rect -142 104 -132 108
rect -82 104 -80 127
rect -78 125 -76 127
rect -70 125 -68 127
rect -63 125 -61 127
rect -66 123 -61 125
rect 17 124 19 126
rect 85 124 87 151
rect 201 143 203 159
rect 226 157 228 159
rect 234 148 236 159
rect 229 144 231 148
rect 234 146 238 148
rect 229 142 234 144
rect 232 140 234 142
rect 236 140 238 146
rect 242 143 244 159
rect 302 143 304 159
rect 327 157 329 159
rect 335 148 337 159
rect 331 144 333 148
rect 335 146 339 148
rect 240 141 244 143
rect 240 140 242 141
rect 201 137 203 139
rect 331 142 335 144
rect 333 140 335 142
rect 337 140 339 146
rect 343 143 345 159
rect 341 141 345 143
rect 341 140 343 141
rect 232 126 234 128
rect -201 103 -199 104
rect -307 89 -305 91
rect -303 73 -301 91
rect -299 73 -297 91
rect -240 70 -238 102
rect -134 102 -132 104
rect -134 96 -132 98
rect -66 96 -64 123
rect 17 122 87 124
rect 158 122 185 124
rect 17 102 19 122
rect 158 120 160 122
rect 183 114 185 122
rect 236 114 238 128
rect 183 112 238 114
rect 158 102 160 108
rect 240 105 242 128
rect 240 103 247 105
rect 4 98 160 102
rect 158 96 160 98
rect -134 94 -64 96
rect -209 89 -207 91
rect -205 73 -203 91
rect -201 73 -199 91
rect 158 88 160 90
rect 4 83 92 87
rect -338 68 -238 70
rect 82 62 84 64
rect 90 62 92 83
rect 98 62 100 87
rect 229 83 231 85
rect 237 83 239 85
rect 245 83 247 103
rect 302 87 304 139
rect 333 126 335 128
rect 337 110 339 128
rect 341 110 343 128
rect 302 85 329 87
rect 204 75 206 77
rect 302 75 304 85
rect 327 83 329 85
rect 335 83 337 85
rect 343 83 345 85
rect 204 65 206 67
rect 229 65 231 67
rect 204 63 231 65
rect 55 54 57 56
rect 128 54 130 56
rect 204 51 206 63
rect 237 56 239 67
rect 233 52 235 56
rect 237 54 241 56
rect 233 50 237 52
rect 235 48 237 50
rect 239 48 241 54
rect 245 51 247 67
rect 302 51 304 67
rect 327 65 329 67
rect 335 56 337 67
rect 331 52 333 56
rect 335 54 339 56
rect 243 49 247 51
rect 243 48 245 49
rect 55 44 57 46
rect 82 44 84 46
rect 55 42 84 44
rect 55 37 57 42
rect 49 33 57 37
rect 90 35 92 46
rect 55 30 57 33
rect 81 31 83 35
rect 90 33 94 35
rect 81 29 90 31
rect 88 27 90 29
rect 92 27 94 33
rect 98 30 100 46
rect 128 36 130 46
rect 120 32 130 36
rect 128 30 130 32
rect 96 28 100 30
rect 96 27 98 28
rect 55 2 57 26
rect 128 24 130 26
rect 88 13 90 15
rect 92 13 94 15
rect 96 13 98 15
rect 204 2 206 47
rect 331 50 335 52
rect 333 48 335 50
rect 337 48 339 54
rect 343 51 345 67
rect 341 49 345 51
rect 341 48 343 49
rect 235 34 237 36
rect 239 18 241 36
rect 243 11 245 36
rect 302 2 304 47
rect 333 34 335 36
rect 337 18 339 36
rect 341 18 343 36
rect 55 0 304 2
<< ndiffusion >>
rect -344 194 -343 198
rect -339 194 -338 198
rect -336 194 -335 198
rect -331 194 -330 198
rect -313 189 -307 195
rect -313 185 -312 189
rect -308 185 -307 189
rect -313 183 -307 185
rect -305 183 -303 195
rect -301 183 -299 195
rect -297 189 -290 195
rect -246 194 -245 198
rect -241 194 -240 198
rect -238 194 -237 198
rect -233 194 -232 198
rect -297 185 -296 189
rect -292 185 -290 189
rect -297 183 -290 185
rect -215 189 -209 195
rect -215 185 -214 189
rect -210 185 -209 189
rect -215 183 -209 185
rect -207 183 -205 195
rect -203 183 -201 195
rect -199 189 -192 195
rect -199 185 -198 189
rect -194 185 -192 189
rect -199 183 -192 185
rect -146 181 -144 185
rect -140 181 -139 185
rect -137 181 -136 185
rect -132 181 -130 185
rect -385 147 -383 151
rect -379 147 -378 151
rect -385 145 -378 147
rect -376 147 -375 151
rect -371 147 -369 151
rect -376 145 -369 147
rect 5 209 7 213
rect 11 209 12 213
rect 14 209 15 213
rect 19 209 21 213
rect 114 170 116 174
rect 120 170 121 174
rect 123 170 124 174
rect 128 170 130 174
rect 51 161 61 167
rect 51 157 56 161
rect 60 157 61 161
rect 51 155 61 157
rect 63 160 69 167
rect 63 156 64 160
rect 68 156 69 160
rect 63 155 69 156
rect 71 155 73 167
rect 75 163 76 167
rect 80 163 81 167
rect 75 155 81 163
rect 83 155 88 167
rect 90 160 95 167
rect 90 156 91 160
rect 90 155 95 156
rect -37 142 -35 146
rect -31 142 -30 146
rect -28 142 -27 146
rect -23 142 -21 146
rect -100 133 -90 139
rect -100 129 -95 133
rect -91 129 -90 133
rect -100 127 -90 129
rect -88 132 -82 139
rect -88 128 -87 132
rect -83 128 -82 132
rect -88 127 -82 128
rect -80 127 -78 139
rect -76 135 -75 139
rect -71 135 -70 139
rect -76 127 -70 135
rect -68 127 -63 139
rect -61 132 -56 139
rect -61 128 -60 132
rect -61 127 -56 128
rect -344 102 -343 106
rect -339 102 -338 106
rect -336 102 -335 106
rect -331 102 -330 106
rect -313 97 -307 103
rect -313 93 -312 97
rect -308 93 -307 97
rect -313 91 -307 93
rect -305 91 -303 103
rect -301 91 -299 103
rect -297 97 -290 103
rect -246 102 -245 106
rect -241 102 -240 106
rect -238 102 -237 106
rect -233 102 -232 106
rect 10 126 12 130
rect 16 126 17 130
rect 19 126 20 130
rect 24 126 26 130
rect 195 139 196 143
rect 200 139 201 143
rect 203 139 204 143
rect 208 139 209 143
rect 226 134 232 140
rect 226 130 227 134
rect 231 130 232 134
rect 226 128 232 130
rect 234 128 236 140
rect 238 128 240 140
rect 242 134 249 140
rect 296 139 297 143
rect 301 139 302 143
rect 304 139 305 143
rect 309 139 310 143
rect 242 130 243 134
rect 247 130 249 134
rect 242 128 249 130
rect -297 93 -296 97
rect -292 93 -290 97
rect -297 91 -290 93
rect -215 97 -209 103
rect -215 93 -214 97
rect -210 93 -209 97
rect -215 91 -209 93
rect -207 91 -205 103
rect -203 91 -201 103
rect -199 97 -192 103
rect -141 98 -139 102
rect -135 98 -134 102
rect -132 98 -131 102
rect -127 98 -125 102
rect -199 93 -198 97
rect -194 93 -192 97
rect -199 91 -192 93
rect 151 92 153 96
rect 157 92 158 96
rect 151 90 158 92
rect 160 92 161 96
rect 165 92 167 96
rect 160 90 167 92
rect 327 134 333 140
rect 327 130 328 134
rect 332 130 333 134
rect 327 128 333 130
rect 335 128 337 140
rect 339 128 341 140
rect 343 134 350 140
rect 343 130 344 134
rect 348 130 350 134
rect 343 128 350 130
rect 198 47 199 51
rect 203 47 204 51
rect 206 47 207 51
rect 211 47 212 51
rect 49 26 50 30
rect 54 26 55 30
rect 57 26 58 30
rect 62 26 63 30
rect 82 21 88 27
rect 82 17 83 21
rect 87 17 88 21
rect 82 15 88 17
rect 90 15 92 27
rect 94 15 96 27
rect 98 21 105 27
rect 122 26 123 30
rect 127 26 128 30
rect 130 26 131 30
rect 135 26 136 30
rect 98 17 99 21
rect 103 17 105 21
rect 98 15 105 17
rect 229 42 235 48
rect 229 38 230 42
rect 234 38 235 42
rect 229 36 235 38
rect 237 36 239 48
rect 241 36 243 48
rect 245 42 252 48
rect 296 47 297 51
rect 301 47 302 51
rect 304 47 305 51
rect 309 47 310 51
rect 245 38 246 42
rect 250 38 252 42
rect 245 36 252 38
rect 327 42 333 48
rect 327 38 328 42
rect 332 38 333 42
rect 327 36 333 38
rect 335 36 337 48
rect 339 36 341 48
rect 343 42 350 48
rect 343 38 344 42
rect 348 38 350 42
rect 343 36 350 38
<< pdiffusion >>
rect -318 229 -313 230
rect -314 225 -313 229
rect -344 218 -343 222
rect -339 218 -338 222
rect -344 214 -338 218
rect -336 218 -335 222
rect -331 218 -330 222
rect -336 214 -330 218
rect -318 214 -313 225
rect -311 229 -305 230
rect -311 225 -310 229
rect -306 225 -305 229
rect -311 214 -305 225
rect -303 220 -297 230
rect -303 216 -302 220
rect -298 216 -297 220
rect -303 214 -297 216
rect -295 229 -290 230
rect -295 225 -294 229
rect -295 214 -290 225
rect -220 229 -215 230
rect -216 225 -215 229
rect -246 218 -245 222
rect -241 218 -240 222
rect -246 214 -240 218
rect -238 218 -237 222
rect -233 218 -232 222
rect -238 214 -232 218
rect -220 214 -215 225
rect -213 229 -207 230
rect -213 225 -212 229
rect -208 225 -207 229
rect -213 214 -207 225
rect -205 220 -199 230
rect -205 216 -204 220
rect -200 216 -199 220
rect -205 214 -199 216
rect -197 229 -192 230
rect -197 225 -196 229
rect -197 214 -192 225
rect -145 205 -144 209
rect -140 205 -139 209
rect -145 201 -139 205
rect -137 205 -136 209
rect -132 205 -131 209
rect -137 201 -131 205
rect -384 171 -383 175
rect -379 171 -378 175
rect -384 163 -378 171
rect -376 171 -375 175
rect -371 171 -370 175
rect -376 163 -370 171
rect -100 173 -95 177
rect -96 169 -95 173
rect -100 153 -95 169
rect -93 172 -87 177
rect -93 168 -92 172
rect -88 168 -87 172
rect -93 153 -87 168
rect -85 165 -79 177
rect -85 161 -84 165
rect -80 161 -79 165
rect -85 153 -79 161
rect -77 157 -71 177
rect -77 153 -76 157
rect -72 153 -71 157
rect -69 165 -63 177
rect -69 161 -68 165
rect -64 161 -63 165
rect -69 153 -63 161
rect -61 172 -56 177
rect -61 168 -60 172
rect 6 233 7 237
rect 11 233 12 237
rect 6 229 12 233
rect 14 233 15 237
rect 19 233 20 237
rect 14 229 20 233
rect 51 201 56 205
rect 55 197 56 201
rect 51 181 56 197
rect 58 200 64 205
rect 58 196 59 200
rect 63 196 64 200
rect 58 181 64 196
rect 66 193 72 205
rect 66 189 67 193
rect 71 189 72 193
rect 66 181 72 189
rect 74 185 80 205
rect 74 181 75 185
rect 79 181 80 185
rect 82 193 88 205
rect 82 189 83 193
rect 87 189 88 193
rect 82 181 88 189
rect 90 200 95 205
rect 90 196 91 200
rect 90 181 95 196
rect 115 194 116 198
rect 120 194 121 198
rect 115 190 121 194
rect 123 194 124 198
rect 128 194 129 198
rect 123 190 129 194
rect -61 153 -56 168
rect -36 166 -35 170
rect -31 166 -30 170
rect -36 162 -30 166
rect -28 166 -27 170
rect -23 166 -22 170
rect -28 162 -22 166
rect -318 137 -313 138
rect -314 133 -313 137
rect -344 126 -343 130
rect -339 126 -338 130
rect -344 122 -338 126
rect -336 126 -335 130
rect -331 126 -330 130
rect -336 122 -330 126
rect -318 122 -313 133
rect -311 137 -305 138
rect -311 133 -310 137
rect -306 133 -305 137
rect -311 122 -305 133
rect -303 128 -297 138
rect -303 124 -302 128
rect -298 124 -297 128
rect -303 122 -297 124
rect -295 137 -290 138
rect -295 133 -294 137
rect -295 122 -290 133
rect -220 137 -215 138
rect -216 133 -215 137
rect -246 126 -245 130
rect -241 126 -240 130
rect -246 122 -240 126
rect -238 126 -237 130
rect -233 126 -232 130
rect -238 122 -232 126
rect -220 122 -215 133
rect -213 137 -207 138
rect -213 133 -212 137
rect -208 133 -207 137
rect -213 122 -207 133
rect -205 128 -199 138
rect -205 124 -204 128
rect -200 124 -199 128
rect -205 122 -199 124
rect -197 137 -192 138
rect -197 133 -196 137
rect -197 122 -192 133
rect 221 174 226 175
rect 225 170 226 174
rect 195 163 196 167
rect 200 163 201 167
rect 195 159 201 163
rect 203 163 204 167
rect 208 163 209 167
rect 203 159 209 163
rect 221 159 226 170
rect 228 174 234 175
rect 228 170 229 174
rect 233 170 234 174
rect 228 159 234 170
rect 236 165 242 175
rect 236 161 237 165
rect 241 161 242 165
rect 236 159 242 161
rect 244 174 249 175
rect 244 170 245 174
rect 244 159 249 170
rect 322 174 327 175
rect 326 170 327 174
rect 296 163 297 167
rect 301 163 302 167
rect 296 159 302 163
rect 304 163 305 167
rect 309 163 310 167
rect 304 159 310 163
rect 322 159 327 170
rect 329 174 335 175
rect 329 170 330 174
rect 334 170 335 174
rect 329 159 335 170
rect 337 165 343 175
rect 337 161 338 165
rect 342 161 343 165
rect 337 159 343 161
rect 345 174 350 175
rect 345 170 346 174
rect 345 159 350 170
rect 11 150 12 154
rect 16 150 17 154
rect 11 146 17 150
rect 19 150 20 154
rect 24 150 25 154
rect 19 146 25 150
rect -140 122 -139 126
rect -135 122 -134 126
rect -140 118 -134 122
rect -132 122 -131 126
rect -127 122 -126 126
rect -132 118 -126 122
rect 152 116 153 120
rect 157 116 158 120
rect 152 108 158 116
rect 160 116 161 120
rect 165 116 166 120
rect 160 108 166 116
rect 224 82 229 83
rect 228 78 229 82
rect 198 71 199 75
rect 203 71 204 75
rect 198 67 204 71
rect 206 71 207 75
rect 211 71 212 75
rect 206 67 212 71
rect 224 67 229 78
rect 231 82 237 83
rect 231 78 232 82
rect 236 78 237 82
rect 231 67 237 78
rect 239 73 245 83
rect 239 69 240 73
rect 244 69 245 73
rect 239 67 245 69
rect 247 82 252 83
rect 247 78 248 82
rect 247 67 252 78
rect 322 82 327 83
rect 326 78 327 82
rect 296 71 297 75
rect 301 71 302 75
rect 296 67 302 71
rect 304 71 305 75
rect 309 71 310 75
rect 304 67 310 71
rect 322 67 327 78
rect 329 82 335 83
rect 329 78 330 82
rect 334 78 335 82
rect 329 67 335 78
rect 337 73 343 83
rect 337 69 338 73
rect 342 69 343 73
rect 337 67 343 69
rect 345 82 350 83
rect 345 78 346 82
rect 345 67 350 78
rect 77 61 82 62
rect 81 57 82 61
rect 49 50 50 54
rect 54 50 55 54
rect 49 46 55 50
rect 57 50 58 54
rect 62 50 63 54
rect 57 46 63 50
rect 77 46 82 57
rect 84 61 90 62
rect 84 57 85 61
rect 89 57 90 61
rect 84 46 90 57
rect 92 52 98 62
rect 92 48 93 52
rect 97 48 98 52
rect 92 46 98 48
rect 100 61 105 62
rect 100 57 101 61
rect 100 46 105 57
rect 122 50 123 54
rect 127 50 128 54
rect 122 46 128 50
rect 130 50 131 54
rect 135 50 136 54
rect 130 46 136 50
<< metal1 >>
rect -30 265 169 269
rect -30 247 -26 265
rect 3 257 23 259
rect 3 253 7 257
rect 11 253 23 257
rect 3 251 23 253
rect -347 242 -281 244
rect -347 238 -343 242
rect -339 238 -318 242
rect -314 238 -294 242
rect -290 238 -281 242
rect -347 236 -281 238
rect -249 242 -183 244
rect -249 238 -245 242
rect -241 238 -220 242
rect -216 238 -196 242
rect -192 238 -183 242
rect -249 236 -183 238
rect 7 237 11 251
rect -343 222 -339 236
rect -318 229 -314 236
rect -306 225 -294 229
rect -245 222 -241 236
rect -220 229 -216 236
rect -148 229 -128 231
rect -208 225 -196 229
rect -148 225 -144 229
rect -140 225 -128 229
rect -148 223 -128 225
rect -335 203 -331 218
rect -302 211 -298 216
rect -302 207 -284 211
rect -288 204 -284 207
rect -335 199 -314 203
rect -288 200 -261 204
rect -335 198 -331 199
rect -387 195 -367 197
rect -387 191 -383 195
rect -379 191 -367 195
rect -387 189 -367 191
rect -383 175 -379 189
rect -343 180 -339 194
rect -288 189 -284 200
rect -292 185 -284 189
rect -312 180 -308 185
rect -347 179 -281 180
rect -347 175 -343 179
rect -339 178 -281 179
rect -339 175 -312 178
rect -347 174 -312 175
rect -308 174 -281 178
rect -347 172 -281 174
rect -375 157 -371 171
rect -265 169 -261 200
rect -237 203 -233 218
rect -204 211 -200 216
rect -204 207 -186 211
rect -190 203 -186 207
rect -144 209 -140 223
rect 15 219 19 233
rect 105 225 143 229
rect -62 215 0 219
rect 15 215 41 219
rect 15 213 19 215
rect -237 199 -215 203
rect -190 199 -166 203
rect -237 198 -233 199
rect -245 180 -241 194
rect -190 189 -186 199
rect -194 185 -186 189
rect -214 180 -210 185
rect -249 179 -183 180
rect -249 175 -245 179
rect -241 178 -183 179
rect -241 175 -214 178
rect -249 174 -214 175
rect -210 174 -183 178
rect -249 172 -183 174
rect -265 165 -209 169
rect -195 165 -176 169
rect -375 153 -358 157
rect -375 151 -371 153
rect -383 133 -379 147
rect -387 132 -367 133
rect -387 128 -383 132
rect -379 128 -367 132
rect -387 125 -367 128
rect -362 77 -358 153
rect -347 150 -281 152
rect -347 146 -343 150
rect -339 146 -318 150
rect -314 146 -294 150
rect -290 146 -281 150
rect -347 144 -281 146
rect -249 150 -183 152
rect -249 146 -245 150
rect -241 146 -220 150
rect -216 146 -196 150
rect -192 146 -183 150
rect -249 144 -183 146
rect -343 130 -339 144
rect -318 137 -314 144
rect -306 133 -294 137
rect -245 130 -241 144
rect -220 137 -216 144
rect -208 133 -196 137
rect -335 111 -331 126
rect -302 119 -298 124
rect -302 115 -284 119
rect -288 112 -284 115
rect -335 107 -313 111
rect -288 108 -263 112
rect -335 106 -331 107
rect -343 88 -339 102
rect -288 97 -284 108
rect -292 93 -284 97
rect -312 88 -308 93
rect -347 87 -281 88
rect -347 83 -343 87
rect -339 86 -281 87
rect -339 83 -312 86
rect -347 82 -312 83
rect -308 82 -281 86
rect -347 80 -281 82
rect -267 77 -263 108
rect -237 111 -233 126
rect -204 119 -200 124
rect -204 115 -186 119
rect -190 112 -186 115
rect -180 112 -176 165
rect -237 107 -215 111
rect -190 108 -176 112
rect -170 108 -166 199
rect -136 191 -132 205
rect -46 197 -8 201
rect -136 187 -110 191
rect -136 185 -132 187
rect -144 167 -140 181
rect -148 166 -128 167
rect -148 162 -144 166
rect -140 162 -128 166
rect -148 159 -128 162
rect -143 146 -123 148
rect -143 142 -139 146
rect -135 142 -123 146
rect -143 140 -123 142
rect -114 144 -110 187
rect -104 189 -60 191
rect -104 185 -100 189
rect -96 185 -60 189
rect -104 183 -60 185
rect -39 190 -19 192
rect -39 186 -35 190
rect -31 186 -19 190
rect -39 184 -19 186
rect -100 173 -96 183
rect -88 168 -60 172
rect -35 170 -31 184
rect -80 161 -68 165
rect -76 148 -72 153
rect -27 152 -23 166
rect -12 152 -8 197
rect 7 195 11 209
rect 3 194 23 195
rect 3 190 7 194
rect 11 190 23 194
rect 3 187 23 190
rect 8 174 28 176
rect 8 170 12 174
rect 16 170 28 174
rect 8 168 28 170
rect 37 172 41 215
rect 47 217 91 219
rect 47 213 51 217
rect 55 213 91 217
rect 47 211 91 213
rect 112 218 132 220
rect 112 214 116 218
rect 120 214 132 218
rect 112 212 132 214
rect 51 201 55 211
rect 63 196 91 200
rect 116 198 120 212
rect 71 189 83 193
rect 75 176 79 181
rect 124 180 128 194
rect 139 180 143 225
rect 75 173 102 176
rect 76 172 102 173
rect 37 168 57 172
rect -27 148 -8 152
rect 12 154 16 168
rect 76 167 80 172
rect 56 150 60 157
rect 68 156 91 160
rect -76 145 -49 148
rect -27 146 -23 148
rect -75 144 -49 145
rect -114 140 -94 144
rect -139 126 -135 140
rect -75 139 -71 144
rect -95 122 -91 129
rect -83 128 -60 132
rect -131 108 -127 122
rect -105 120 -61 122
rect -105 116 -95 120
rect -91 116 -61 120
rect -105 114 -61 116
rect -237 106 -233 107
rect -245 88 -241 102
rect -190 97 -186 108
rect -194 93 -186 97
rect -170 104 -146 108
rect -131 104 -86 108
rect -214 88 -210 93
rect -249 87 -183 88
rect -249 83 -245 87
rect -241 86 -183 87
rect -241 83 -214 86
rect -249 82 -214 83
rect -210 82 -183 86
rect -249 80 -183 82
rect -170 77 -166 104
rect -131 102 -127 104
rect -53 102 -49 144
rect -35 128 -31 142
rect 20 136 24 150
rect 46 148 90 150
rect 46 144 56 148
rect 60 144 90 148
rect 46 142 90 144
rect 20 132 65 136
rect 20 130 24 132
rect -39 127 -19 128
rect -39 123 -35 127
rect -31 123 -19 127
rect -39 120 -19 123
rect 12 112 16 126
rect 98 121 102 172
rect 109 162 113 176
rect 124 176 143 180
rect 165 196 169 265
rect 165 192 376 196
rect 124 174 128 176
rect 105 159 113 162
rect 105 144 109 159
rect 116 156 120 170
rect 112 155 132 156
rect 112 151 116 155
rect 120 151 132 155
rect 165 154 169 192
rect 192 187 258 189
rect 192 183 196 187
rect 200 183 221 187
rect 225 183 245 187
rect 249 183 258 187
rect 192 181 258 183
rect 293 187 359 189
rect 293 183 297 187
rect 301 183 322 187
rect 326 183 346 187
rect 350 183 359 187
rect 293 181 359 183
rect 196 167 200 181
rect 221 174 225 181
rect 233 170 245 174
rect 297 167 301 181
rect 322 174 326 181
rect 334 170 346 174
rect 112 148 132 151
rect 138 150 169 154
rect 138 144 142 150
rect 105 140 142 144
rect 204 148 208 163
rect 237 156 241 161
rect 237 152 255 156
rect 251 149 255 152
rect 204 144 225 148
rect 251 145 281 149
rect 204 143 208 144
rect 149 140 169 142
rect 149 136 153 140
rect 157 136 169 140
rect 149 134 169 136
rect 98 117 104 121
rect 8 111 28 112
rect 8 107 12 111
rect 16 107 28 111
rect 8 104 28 107
rect -53 98 0 102
rect -139 84 -135 98
rect 100 87 104 117
rect 153 120 157 134
rect 196 125 200 139
rect 251 134 255 145
rect 247 130 255 134
rect 227 125 231 130
rect 192 124 258 125
rect 192 120 196 124
rect 200 123 258 124
rect 200 120 227 123
rect 192 119 227 120
rect 231 119 258 123
rect 192 117 258 119
rect 161 102 165 116
rect 277 114 281 145
rect 305 148 309 163
rect 338 156 342 161
rect 338 152 356 156
rect 352 148 356 152
rect 372 148 376 192
rect 305 144 327 148
rect 352 144 380 148
rect 305 143 309 144
rect 297 125 301 139
rect 352 134 356 144
rect 348 130 356 134
rect 328 125 332 130
rect 293 124 359 125
rect 293 120 297 124
rect 301 123 359 124
rect 301 120 328 123
rect 293 119 328 120
rect 332 119 359 123
rect 293 117 359 119
rect 277 110 333 114
rect 347 110 366 114
rect 161 98 184 102
rect 161 96 165 98
rect -362 73 -307 77
rect -267 73 -209 77
rect -195 73 -166 77
rect -143 83 -123 84
rect -143 79 -139 83
rect -135 79 -123 83
rect -143 76 -123 79
rect -23 83 0 87
rect -297 66 -293 73
rect -23 66 -19 83
rect 153 78 157 92
rect 149 77 169 78
rect 46 74 139 76
rect 46 70 50 74
rect 54 70 77 74
rect 81 70 101 74
rect 105 70 123 74
rect 127 70 139 74
rect 149 73 153 77
rect 157 73 169 77
rect 149 70 169 73
rect 46 68 139 70
rect -297 62 -19 66
rect 50 54 54 68
rect 77 61 81 68
rect 89 57 101 61
rect 123 54 127 68
rect 58 35 62 50
rect 93 43 97 48
rect 93 39 111 43
rect 107 36 111 39
rect 131 36 135 50
rect 58 31 77 35
rect 107 32 116 36
rect 107 31 120 32
rect 131 32 156 36
rect 58 30 62 31
rect 50 12 54 26
rect 107 21 111 31
rect 131 30 135 32
rect 103 17 111 21
rect 83 12 87 17
rect 123 12 127 26
rect 152 15 156 32
rect 180 22 184 98
rect 195 95 261 97
rect 195 91 199 95
rect 203 91 224 95
rect 228 91 248 95
rect 252 91 261 95
rect 195 89 261 91
rect 293 95 359 97
rect 293 91 297 95
rect 301 91 322 95
rect 326 91 346 95
rect 350 91 359 95
rect 293 89 359 91
rect 199 75 203 89
rect 224 82 228 89
rect 236 78 248 82
rect 297 75 301 89
rect 322 82 326 89
rect 334 78 346 82
rect 207 56 211 71
rect 240 64 244 69
rect 240 60 258 64
rect 254 57 258 60
rect 207 52 229 56
rect 254 53 279 57
rect 207 51 211 52
rect 199 33 203 47
rect 254 42 258 53
rect 250 38 258 42
rect 230 33 234 38
rect 195 32 261 33
rect 195 28 199 32
rect 203 31 261 32
rect 203 28 230 31
rect 195 27 230 28
rect 234 27 261 31
rect 195 25 261 27
rect 275 22 279 53
rect 305 56 309 71
rect 338 64 342 69
rect 338 60 356 64
rect 352 57 356 60
rect 362 57 366 110
rect 305 52 327 56
rect 352 53 366 57
rect 305 51 309 52
rect 297 33 301 47
rect 352 42 356 53
rect 348 38 356 42
rect 328 33 332 38
rect 293 32 359 33
rect 293 28 297 32
rect 301 31 359 32
rect 301 28 328 31
rect 293 27 328 28
rect 332 27 359 31
rect 293 25 359 27
rect 372 22 376 144
rect 180 18 235 22
rect 275 18 333 22
rect 347 18 376 22
rect 46 11 139 12
rect 152 11 239 15
rect 46 7 50 11
rect 54 10 123 11
rect 54 7 83 10
rect 46 6 83 7
rect 87 7 123 10
rect 127 7 139 11
rect 87 6 139 7
rect 46 4 139 6
<< ntransistor >>
rect -338 194 -336 198
rect -307 183 -305 195
rect -303 183 -301 195
rect -299 183 -297 195
rect -240 194 -238 198
rect -209 183 -207 195
rect -205 183 -203 195
rect -201 183 -199 195
rect -139 181 -137 185
rect -378 145 -376 151
rect 12 209 14 213
rect 121 170 123 174
rect 61 155 63 167
rect 69 155 71 167
rect 73 155 75 167
rect 81 155 83 167
rect 88 155 90 167
rect -30 142 -28 146
rect -90 127 -88 139
rect -82 127 -80 139
rect -78 127 -76 139
rect -70 127 -68 139
rect -63 127 -61 139
rect -338 102 -336 106
rect -307 91 -305 103
rect -303 91 -301 103
rect -299 91 -297 103
rect -240 102 -238 106
rect 17 126 19 130
rect 201 139 203 143
rect 232 128 234 140
rect 236 128 238 140
rect 240 128 242 140
rect 302 139 304 143
rect -209 91 -207 103
rect -205 91 -203 103
rect -201 91 -199 103
rect -134 98 -132 102
rect 158 90 160 96
rect 333 128 335 140
rect 337 128 339 140
rect 341 128 343 140
rect 204 47 206 51
rect 55 26 57 30
rect 88 15 90 27
rect 92 15 94 27
rect 96 15 98 27
rect 128 26 130 30
rect 235 36 237 48
rect 239 36 241 48
rect 243 36 245 48
rect 302 47 304 51
rect 333 36 335 48
rect 337 36 339 48
rect 341 36 343 48
<< ptransistor >>
rect -338 214 -336 222
rect -313 214 -311 230
rect -305 214 -303 230
rect -297 214 -295 230
rect -240 214 -238 222
rect -215 214 -213 230
rect -207 214 -205 230
rect -199 214 -197 230
rect -139 201 -137 209
rect -378 163 -376 175
rect -95 153 -93 177
rect -87 153 -85 177
rect -79 153 -77 177
rect -71 153 -69 177
rect -63 153 -61 177
rect 12 229 14 237
rect 56 181 58 205
rect 64 181 66 205
rect 72 181 74 205
rect 80 181 82 205
rect 88 181 90 205
rect 121 190 123 198
rect -30 162 -28 170
rect -338 122 -336 130
rect -313 122 -311 138
rect -305 122 -303 138
rect -297 122 -295 138
rect -240 122 -238 130
rect -215 122 -213 138
rect -207 122 -205 138
rect -199 122 -197 138
rect 201 159 203 167
rect 226 159 228 175
rect 234 159 236 175
rect 242 159 244 175
rect 302 159 304 167
rect 327 159 329 175
rect 335 159 337 175
rect 343 159 345 175
rect 17 146 19 154
rect -134 118 -132 126
rect 158 108 160 120
rect 204 67 206 75
rect 229 67 231 83
rect 237 67 239 83
rect 245 67 247 83
rect 302 67 304 75
rect 327 67 329 83
rect 335 67 337 83
rect 343 67 345 83
rect 55 46 57 54
rect 82 46 84 62
rect 90 46 92 62
rect 98 46 100 62
rect 128 46 130 54
<< polycontact >>
rect -30 243 -26 247
rect -314 199 -310 203
rect -215 199 -211 203
rect -66 215 -62 219
rect -303 158 -299 162
rect -50 197 -46 201
rect -209 165 -205 169
rect -199 165 -195 169
rect -383 154 -379 158
rect 0 215 4 219
rect 101 225 105 229
rect -94 140 -90 144
rect 57 168 61 172
rect 109 176 113 180
rect -42 148 -38 152
rect 65 132 69 136
rect -313 107 -309 111
rect -215 107 -211 111
rect -146 104 -142 108
rect -86 104 -82 108
rect 225 144 229 148
rect 327 144 331 148
rect -307 73 -303 77
rect -297 73 -293 77
rect 0 98 4 102
rect -209 73 -205 77
rect 0 83 4 87
rect -199 73 -195 77
rect 100 83 104 87
rect 333 110 337 114
rect 343 110 347 114
rect 229 52 233 56
rect 327 52 331 56
rect 45 33 49 37
rect 77 31 81 35
rect 116 32 120 36
rect 235 18 239 22
rect 239 11 243 15
rect 333 18 337 22
rect 343 18 347 22
<< ndcontact >>
rect -343 194 -339 198
rect -335 194 -331 198
rect -312 185 -308 189
rect -245 194 -241 198
rect -237 194 -233 198
rect -296 185 -292 189
rect -214 185 -210 189
rect -198 185 -194 189
rect -144 181 -140 185
rect -136 181 -132 185
rect -383 147 -379 151
rect -375 147 -371 151
rect 7 209 11 213
rect 15 209 19 213
rect 116 170 120 174
rect 124 170 128 174
rect 56 157 60 161
rect 64 156 68 160
rect 76 163 80 167
rect 91 156 95 160
rect -35 142 -31 146
rect -27 142 -23 146
rect -95 129 -91 133
rect -87 128 -83 132
rect -75 135 -71 139
rect -60 128 -56 132
rect -343 102 -339 106
rect -335 102 -331 106
rect -312 93 -308 97
rect -245 102 -241 106
rect -237 102 -233 106
rect 12 126 16 130
rect 20 126 24 130
rect 196 139 200 143
rect 204 139 208 143
rect 227 130 231 134
rect 297 139 301 143
rect 305 139 309 143
rect 243 130 247 134
rect -296 93 -292 97
rect -214 93 -210 97
rect -139 98 -135 102
rect -131 98 -127 102
rect -198 93 -194 97
rect 153 92 157 96
rect 161 92 165 96
rect 328 130 332 134
rect 344 130 348 134
rect 199 47 203 51
rect 207 47 211 51
rect 50 26 54 30
rect 58 26 62 30
rect 83 17 87 21
rect 123 26 127 30
rect 131 26 135 30
rect 99 17 103 21
rect 230 38 234 42
rect 297 47 301 51
rect 305 47 309 51
rect 246 38 250 42
rect 328 38 332 42
rect 344 38 348 42
<< pdcontact >>
rect -318 225 -314 229
rect -343 218 -339 222
rect -335 218 -331 222
rect -310 225 -306 229
rect -302 216 -298 220
rect -294 225 -290 229
rect -220 225 -216 229
rect -245 218 -241 222
rect -237 218 -233 222
rect -212 225 -208 229
rect -204 216 -200 220
rect -196 225 -192 229
rect -144 205 -140 209
rect -136 205 -132 209
rect -383 171 -379 175
rect -375 171 -371 175
rect -100 169 -96 173
rect -92 168 -88 172
rect -84 161 -80 165
rect -76 153 -72 157
rect -68 161 -64 165
rect -60 168 -56 172
rect 7 233 11 237
rect 15 233 19 237
rect 51 197 55 201
rect 59 196 63 200
rect 67 189 71 193
rect 75 181 79 185
rect 83 189 87 193
rect 91 196 95 200
rect 116 194 120 198
rect 124 194 128 198
rect -35 166 -31 170
rect -27 166 -23 170
rect -318 133 -314 137
rect -343 126 -339 130
rect -335 126 -331 130
rect -310 133 -306 137
rect -302 124 -298 128
rect -294 133 -290 137
rect -220 133 -216 137
rect -245 126 -241 130
rect -237 126 -233 130
rect -212 133 -208 137
rect -204 124 -200 128
rect -196 133 -192 137
rect 221 170 225 174
rect 196 163 200 167
rect 204 163 208 167
rect 229 170 233 174
rect 237 161 241 165
rect 245 170 249 174
rect 322 170 326 174
rect 297 163 301 167
rect 305 163 309 167
rect 330 170 334 174
rect 338 161 342 165
rect 346 170 350 174
rect 12 150 16 154
rect 20 150 24 154
rect -139 122 -135 126
rect -131 122 -127 126
rect 153 116 157 120
rect 161 116 165 120
rect 224 78 228 82
rect 199 71 203 75
rect 207 71 211 75
rect 232 78 236 82
rect 240 69 244 73
rect 248 78 252 82
rect 322 78 326 82
rect 297 71 301 75
rect 305 71 309 75
rect 330 78 334 82
rect 338 69 342 73
rect 346 78 350 82
rect 77 57 81 61
rect 50 50 54 54
rect 58 50 62 54
rect 85 57 89 61
rect 93 48 97 52
rect 101 57 105 61
rect 123 50 127 54
rect 131 50 135 54
<< psubstratepcontact >>
rect -343 175 -339 179
rect -312 174 -308 178
rect -245 175 -241 179
rect -214 174 -210 178
rect -144 162 -140 166
rect 7 190 11 194
rect -383 128 -379 132
rect 56 144 60 148
rect 116 151 120 155
rect -343 83 -339 87
rect -95 116 -91 120
rect -35 123 -31 127
rect -312 82 -308 86
rect -245 83 -241 87
rect 12 107 16 111
rect 196 120 200 124
rect 227 119 231 123
rect 297 120 301 124
rect -214 82 -210 86
rect -139 79 -135 83
rect 328 119 332 123
rect 153 73 157 77
rect 50 7 54 11
rect 199 28 203 32
rect 83 6 87 10
rect 123 7 127 11
rect 230 27 234 31
rect 297 28 301 32
rect 328 27 332 31
<< nsubstratencontact >>
rect 7 253 11 257
rect -383 191 -379 195
rect -343 238 -339 242
rect -318 238 -314 242
rect -294 238 -290 242
rect -245 238 -241 242
rect -220 238 -216 242
rect -196 238 -192 242
rect -144 225 -140 229
rect -100 185 -96 189
rect -35 186 -31 190
rect -343 146 -339 150
rect -318 146 -314 150
rect -294 146 -290 150
rect -245 146 -241 150
rect 51 213 55 217
rect 116 214 120 218
rect 12 170 16 174
rect -220 146 -216 150
rect -196 146 -192 150
rect -139 142 -135 146
rect 196 183 200 187
rect 221 183 225 187
rect 245 183 249 187
rect 297 183 301 187
rect 322 183 326 187
rect 346 183 350 187
rect 153 136 157 140
rect 199 91 203 95
rect 224 91 228 95
rect 50 70 54 74
rect 77 70 81 74
rect 248 91 252 95
rect 297 91 301 95
rect 322 91 326 95
rect 346 91 350 95
rect 101 70 105 74
rect 123 70 127 74
<< labels >>
rlabel nwell 192 181 258 189 1 vdd_1
rlabel nwell 293 181 359 189 1 vdd_2
rlabel nwell 293 89 359 97 1 vdd_4
rlabel nwell 195 89 261 97 1 vdd_3
rlabel metal1 192 117 258 125 5 vss_1
rlabel metal1 293 117 359 125 5 vss_2
rlabel metal1 293 25 359 33 5 vss_4
rlabel metal1 195 25 261 33 5 vss_3
rlabel polycontact 239 11 243 15 5 gated_clk
rlabel metal1 149 70 169 78 5 vss_5
rlabel nwell 149 134 169 142 1 vdd_5
rlabel nwell 46 68 139 76 1 vdd_10
rlabel metal1 46 4 139 12 5 vss_10
rlabel polycontact 0 215 4 219 5 sleep
rlabel nwell 3 251 23 259 1 vdd_6
rlabel metal1 3 187 23 195 5 vss_6
rlabel nwell 8 168 28 176 1 vdd_7
rlabel metal1 8 104 28 112 5 vss_7
rlabel metal1 47 211 91 219 1 vdd_8
rlabel metal1 46 142 90 150 5 vss_8
rlabel nwell 112 212 132 220 1 vdd_9
rlabel metal1 112 148 132 156 5 vss_9
rlabel polycontact 0 83 4 87 5 clk
rlabel nwell -387 189 -367 197 1 vdd_11
rlabel metal1 -387 125 -367 133 5 vss_11
rlabel nwell -347 236 -281 244 1 vdd_12
rlabel nwell -249 236 -183 244 1 vdd_13
rlabel nwell -347 144 -281 152 1 vdd_14
rlabel nwell -249 144 -183 152 1 vdd_15
rlabel metal1 -347 172 -281 180 5 vss_12
rlabel metal1 -249 172 -183 180 5 vss_13
rlabel metal1 -347 80 -281 88 5 vss_14
rlabel metal1 -249 80 -183 88 5 vss_15
rlabel nwell -148 223 -128 231 1 vdd_16
rlabel nwell -143 140 -123 148 1 vdd_17
rlabel metal1 -104 183 -60 191 1 vdd_18
rlabel nwell -39 184 -19 192 1 vdd_19
rlabel metal1 -148 159 -128 167 5 vss_16
rlabel metal1 -143 76 -123 84 5 vss_17
rlabel metal1 -39 120 -19 128 5 vss_19
rlabel metal1 -105 114 -61 122 5 vss_18
rlabel metal1 376 144 380 148 3 out_1
rlabel polycontact -146 104 -142 108 5 out_0
rlabel polycontact -383 154 -379 158 7 d
rlabel polycontact 0 98 4 102 5 d2
rlabel polycontact 100 83 104 87 3 desn
<< end >>
