magic
tech scmos
timestamp 1679571716
<< nwell >>
rect 109 19 178 50
rect 207 19 276 50
rect 109 12 136 19
rect 207 12 234 19
rect 69 -35 96 6
rect 109 -73 178 -42
rect 207 -73 276 -42
rect 109 -80 136 -73
rect 207 -80 234 -73
<< polysilicon >>
rect 121 40 221 42
rect 121 28 123 40
rect 146 36 148 40
rect 219 38 246 40
rect 154 36 156 38
rect 162 36 164 38
rect 219 28 221 38
rect 244 36 246 38
rect 252 36 254 38
rect 260 36 262 38
rect 121 10 123 20
rect 146 18 148 20
rect 113 6 123 10
rect 154 9 156 20
rect 121 4 123 6
rect 149 5 151 9
rect 154 7 158 9
rect 149 3 154 5
rect 152 1 154 3
rect 156 1 158 7
rect 162 4 164 20
rect 219 4 221 20
rect 244 18 246 20
rect 252 9 254 20
rect 248 5 250 9
rect 252 7 256 9
rect 160 2 164 4
rect 160 1 162 2
rect 121 -2 123 0
rect 248 3 252 5
rect 250 1 252 3
rect 254 1 256 7
rect 260 4 262 20
rect 258 2 262 4
rect 258 1 260 2
rect 152 -13 154 -11
rect 81 -17 105 -15
rect 81 -19 83 -17
rect 103 -25 105 -17
rect 156 -25 158 -11
rect 103 -27 158 -25
rect 81 -37 83 -31
rect 160 -34 162 -11
rect 160 -36 164 -34
rect 73 -41 83 -37
rect 81 -43 83 -41
rect 81 -52 83 -49
rect 146 -56 148 -54
rect 154 -56 156 -54
rect 162 -56 164 -36
rect 219 -52 221 0
rect 250 -13 252 -11
rect 254 -29 256 -11
rect 258 -29 260 -11
rect 219 -54 246 -52
rect 121 -64 123 -62
rect 219 -64 221 -54
rect 244 -56 246 -54
rect 252 -56 254 -54
rect 260 -56 262 -54
rect 121 -74 123 -72
rect 146 -74 148 -72
rect 121 -76 148 -74
rect 121 -88 123 -76
rect 154 -83 156 -72
rect 150 -87 152 -83
rect 154 -85 158 -83
rect 150 -89 154 -87
rect 152 -91 154 -89
rect 156 -91 158 -85
rect 162 -88 164 -72
rect 219 -88 221 -72
rect 244 -74 246 -72
rect 252 -83 254 -72
rect 248 -87 250 -83
rect 252 -85 256 -83
rect 160 -90 164 -88
rect 160 -91 162 -90
rect 121 -124 123 -92
rect 248 -89 252 -87
rect 250 -91 252 -89
rect 254 -91 256 -85
rect 260 -88 262 -72
rect 258 -90 262 -88
rect 258 -91 260 -90
rect 152 -105 154 -103
rect 156 -121 158 -103
rect 160 -116 162 -103
rect 219 -124 221 -92
rect 250 -105 252 -103
rect 254 -121 256 -103
rect 258 -121 260 -103
rect 121 -126 221 -124
<< ndiffusion >>
rect 115 0 116 4
rect 120 0 121 4
rect 123 0 124 4
rect 128 0 129 4
rect 146 -5 152 1
rect 146 -9 147 -5
rect 151 -9 152 -5
rect 146 -11 152 -9
rect 154 -11 156 1
rect 158 -11 160 1
rect 162 -5 169 1
rect 213 0 214 4
rect 218 0 219 4
rect 221 0 222 4
rect 226 0 227 4
rect 162 -9 163 -5
rect 167 -9 169 -5
rect 162 -11 169 -9
rect 74 -47 76 -43
rect 80 -47 81 -43
rect 74 -49 81 -47
rect 83 -47 84 -43
rect 88 -47 90 -43
rect 83 -49 90 -47
rect 244 -5 250 1
rect 244 -9 245 -5
rect 249 -9 250 -5
rect 244 -11 250 -9
rect 252 -11 254 1
rect 256 -11 258 1
rect 260 -5 267 1
rect 260 -9 261 -5
rect 265 -9 267 -5
rect 260 -11 267 -9
rect 115 -92 116 -88
rect 120 -92 121 -88
rect 123 -92 124 -88
rect 128 -92 129 -88
rect 146 -97 152 -91
rect 146 -101 147 -97
rect 151 -101 152 -97
rect 146 -103 152 -101
rect 154 -103 156 -91
rect 158 -103 160 -91
rect 162 -97 169 -91
rect 213 -92 214 -88
rect 218 -92 219 -88
rect 221 -92 222 -88
rect 226 -92 227 -88
rect 162 -101 163 -97
rect 167 -101 169 -97
rect 162 -103 169 -101
rect 244 -97 250 -91
rect 244 -101 245 -97
rect 249 -101 250 -97
rect 244 -103 250 -101
rect 252 -103 254 -91
rect 256 -103 258 -91
rect 260 -97 267 -91
rect 260 -101 261 -97
rect 265 -101 267 -97
rect 260 -103 267 -101
<< pdiffusion >>
rect 141 35 146 36
rect 145 31 146 35
rect 115 24 116 28
rect 120 24 121 28
rect 115 20 121 24
rect 123 24 124 28
rect 128 24 129 28
rect 123 20 129 24
rect 141 20 146 31
rect 148 35 154 36
rect 148 31 149 35
rect 153 31 154 35
rect 148 20 154 31
rect 156 26 162 36
rect 156 22 157 26
rect 161 22 162 26
rect 156 20 162 22
rect 164 35 169 36
rect 164 31 165 35
rect 164 20 169 31
rect 239 35 244 36
rect 243 31 244 35
rect 213 24 214 28
rect 218 24 219 28
rect 213 20 219 24
rect 221 24 222 28
rect 226 24 227 28
rect 221 20 227 24
rect 239 20 244 31
rect 246 35 252 36
rect 246 31 247 35
rect 251 31 252 35
rect 246 20 252 31
rect 254 26 260 36
rect 254 22 255 26
rect 259 22 260 26
rect 254 20 260 22
rect 262 35 267 36
rect 262 31 263 35
rect 262 20 267 31
rect 75 -23 76 -19
rect 80 -23 81 -19
rect 75 -31 81 -23
rect 83 -23 84 -19
rect 88 -23 89 -19
rect 83 -31 89 -23
rect 141 -57 146 -56
rect 145 -61 146 -57
rect 115 -68 116 -64
rect 120 -68 121 -64
rect 115 -72 121 -68
rect 123 -68 124 -64
rect 128 -68 129 -64
rect 123 -72 129 -68
rect 141 -72 146 -61
rect 148 -57 154 -56
rect 148 -61 149 -57
rect 153 -61 154 -57
rect 148 -72 154 -61
rect 156 -66 162 -56
rect 156 -70 157 -66
rect 161 -70 162 -66
rect 156 -72 162 -70
rect 164 -57 169 -56
rect 164 -61 165 -57
rect 164 -72 169 -61
rect 239 -57 244 -56
rect 243 -61 244 -57
rect 213 -68 214 -64
rect 218 -68 219 -64
rect 213 -72 219 -68
rect 221 -68 222 -64
rect 226 -68 227 -64
rect 221 -72 227 -68
rect 239 -72 244 -61
rect 246 -57 252 -56
rect 246 -61 247 -57
rect 251 -61 252 -57
rect 246 -72 252 -61
rect 254 -66 260 -56
rect 254 -70 255 -66
rect 259 -70 260 -66
rect 254 -72 260 -70
rect 262 -57 267 -56
rect 262 -61 263 -57
rect 262 -72 267 -61
<< metal1 >>
rect 112 48 178 50
rect 112 44 116 48
rect 120 44 141 48
rect 145 44 165 48
rect 169 44 178 48
rect 112 42 178 44
rect 210 48 276 50
rect 210 44 214 48
rect 218 44 239 48
rect 243 44 263 48
rect 267 44 276 48
rect 210 42 276 44
rect 116 28 120 42
rect 141 35 145 42
rect 153 31 165 35
rect 214 28 218 42
rect 239 35 243 42
rect 251 31 263 35
rect 124 9 128 24
rect 157 17 161 22
rect 157 13 175 17
rect 171 10 175 13
rect 124 5 145 9
rect 171 6 198 10
rect 124 4 128 5
rect 72 1 92 3
rect 72 -3 76 1
rect 80 -3 92 1
rect 72 -5 92 -3
rect 76 -19 80 -5
rect 116 -14 120 0
rect 171 -5 175 6
rect 167 -9 175 -5
rect 147 -14 151 -9
rect 112 -15 178 -14
rect 112 -19 116 -15
rect 120 -16 178 -15
rect 120 -19 147 -16
rect 112 -20 147 -19
rect 151 -20 178 -16
rect 112 -22 178 -20
rect 84 -37 88 -23
rect 194 -25 198 6
rect 222 9 226 24
rect 255 17 259 22
rect 255 13 273 17
rect 269 9 273 13
rect 222 5 244 9
rect 269 5 297 9
rect 222 4 226 5
rect 214 -14 218 0
rect 269 -5 273 5
rect 265 -9 273 -5
rect 245 -14 249 -9
rect 210 -15 276 -14
rect 210 -19 214 -15
rect 218 -16 276 -15
rect 218 -19 245 -16
rect 210 -20 245 -19
rect 249 -20 276 -16
rect 210 -22 276 -20
rect 194 -29 250 -25
rect 264 -29 283 -25
rect 84 -41 101 -37
rect 84 -43 88 -41
rect 76 -61 80 -47
rect 72 -62 92 -61
rect 72 -66 76 -62
rect 80 -66 92 -62
rect 72 -69 92 -66
rect 97 -117 101 -41
rect 112 -44 178 -42
rect 112 -48 116 -44
rect 120 -48 141 -44
rect 145 -48 165 -44
rect 169 -48 178 -44
rect 112 -50 178 -48
rect 210 -44 276 -42
rect 210 -48 214 -44
rect 218 -48 239 -44
rect 243 -48 263 -44
rect 267 -48 276 -44
rect 210 -50 276 -48
rect 116 -64 120 -50
rect 141 -57 145 -50
rect 153 -61 165 -57
rect 214 -64 218 -50
rect 239 -57 243 -50
rect 251 -61 263 -57
rect 124 -83 128 -68
rect 157 -75 161 -70
rect 157 -79 175 -75
rect 171 -82 175 -79
rect 124 -87 146 -83
rect 171 -86 196 -82
rect 124 -88 128 -87
rect 116 -106 120 -92
rect 171 -97 175 -86
rect 167 -101 175 -97
rect 147 -106 151 -101
rect 112 -107 178 -106
rect 112 -111 116 -107
rect 120 -108 178 -107
rect 120 -111 147 -108
rect 112 -112 147 -111
rect 151 -112 178 -108
rect 112 -114 178 -112
rect 192 -117 196 -86
rect 222 -83 226 -68
rect 255 -75 259 -70
rect 255 -79 273 -75
rect 269 -82 273 -79
rect 279 -82 283 -29
rect 222 -87 244 -83
rect 269 -86 283 -82
rect 222 -88 226 -87
rect 214 -106 218 -92
rect 269 -97 273 -86
rect 265 -101 273 -97
rect 245 -106 249 -101
rect 210 -107 276 -106
rect 210 -111 214 -107
rect 218 -108 276 -107
rect 218 -111 245 -108
rect 210 -112 245 -111
rect 249 -112 276 -108
rect 210 -114 276 -112
rect 289 -117 293 5
rect 97 -121 152 -117
rect 192 -121 250 -117
rect 264 -121 293 -117
<< ntransistor >>
rect 121 0 123 4
rect 152 -11 154 1
rect 156 -11 158 1
rect 160 -11 162 1
rect 219 0 221 4
rect 81 -49 83 -43
rect 250 -11 252 1
rect 254 -11 256 1
rect 258 -11 260 1
rect 121 -92 123 -88
rect 152 -103 154 -91
rect 156 -103 158 -91
rect 160 -103 162 -91
rect 219 -92 221 -88
rect 250 -103 252 -91
rect 254 -103 256 -91
rect 258 -103 260 -91
<< ptransistor >>
rect 121 20 123 28
rect 146 20 148 36
rect 154 20 156 36
rect 162 20 164 36
rect 219 20 221 28
rect 244 20 246 36
rect 252 20 254 36
rect 260 20 262 36
rect 81 -31 83 -19
rect 121 -72 123 -64
rect 146 -72 148 -56
rect 154 -72 156 -56
rect 162 -72 164 -56
rect 219 -72 221 -64
rect 244 -72 246 -56
rect 252 -72 254 -56
rect 260 -72 262 -56
<< polycontact >>
rect 109 6 113 10
rect 145 5 149 9
rect 244 5 248 9
rect 156 -36 160 -32
rect 69 -41 73 -37
rect 250 -29 254 -25
rect 260 -29 264 -25
rect 146 -87 150 -83
rect 244 -87 248 -83
rect 152 -121 156 -117
rect 250 -121 254 -117
rect 260 -121 264 -117
<< ndcontact >>
rect 116 0 120 4
rect 124 0 128 4
rect 147 -9 151 -5
rect 214 0 218 4
rect 222 0 226 4
rect 163 -9 167 -5
rect 76 -47 80 -43
rect 84 -47 88 -43
rect 245 -9 249 -5
rect 261 -9 265 -5
rect 116 -92 120 -88
rect 124 -92 128 -88
rect 147 -101 151 -97
rect 214 -92 218 -88
rect 222 -92 226 -88
rect 163 -101 167 -97
rect 245 -101 249 -97
rect 261 -101 265 -97
<< pdcontact >>
rect 141 31 145 35
rect 116 24 120 28
rect 124 24 128 28
rect 149 31 153 35
rect 157 22 161 26
rect 165 31 169 35
rect 239 31 243 35
rect 214 24 218 28
rect 222 24 226 28
rect 247 31 251 35
rect 255 22 259 26
rect 263 31 267 35
rect 76 -23 80 -19
rect 84 -23 88 -19
rect 141 -61 145 -57
rect 116 -68 120 -64
rect 124 -68 128 -64
rect 149 -61 153 -57
rect 157 -70 161 -66
rect 165 -61 169 -57
rect 239 -61 243 -57
rect 214 -68 218 -64
rect 222 -68 226 -64
rect 247 -61 251 -57
rect 255 -70 259 -66
rect 263 -61 267 -57
<< psubstratepcontact >>
rect 116 -19 120 -15
rect 147 -20 151 -16
rect 214 -19 218 -15
rect 245 -20 249 -16
rect 76 -66 80 -62
rect 116 -111 120 -107
rect 147 -112 151 -108
rect 214 -111 218 -107
rect 245 -112 249 -108
<< nsubstratencontact >>
rect 116 44 120 48
rect 141 44 145 48
rect 165 44 169 48
rect 214 44 218 48
rect 239 44 243 48
rect 263 44 267 48
rect 76 -3 80 1
rect 116 -48 120 -44
rect 141 -48 145 -44
rect 165 -48 169 -44
rect 214 -48 218 -44
rect 239 -48 243 -44
rect 263 -48 267 -44
<< labels >>
rlabel nwell 210 42 276 50 1 vdd_2
rlabel nwell 210 -50 276 -42 1 vdd_4
rlabel metal1 210 -22 276 -14 5 vss_2
rlabel metal1 210 -114 276 -106 5 vss_4
rlabel metal1 112 -114 178 -106 5 vss_3
rlabel metal1 293 5 297 9 3 out
rlabel nwell 112 -50 178 -42 1 vdd_3
rlabel nwell 112 42 178 50 1 vdd_1
rlabel polycontact 109 6 113 10 5 slp
rlabel metal1 112 -22 178 -14 5 vss_1
rlabel polycontact 156 -36 160 -32 5 clock
rlabel metal1 72 -69 92 -61 5 vss
rlabel nwell 72 -5 92 3 1 vdd
rlabel metal1 88 -41 91 -37 5 d_n
rlabel polycontact 69 -41 73 -37 5 d
rlabel metal1 279 -86 283 -82 5 out_n
<< end >>
